-- $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/vhdsclibs/data/simprims/stan/SMODEL/X_MCB.vhd,v 1.11 2010/02/04 21:02:42 vandanad Exp $
-------------------------------------------------------
--  Copyright (c) 2008 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version : 11.1
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : X_MCB.vhd
-- \   \  /  \      
--  \__ \/\__ \                   
--                                 
--  Generated by    : /home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/write_vhdl.pl
--  Revision: 1.0
--  518974 - X_MCB.vhd - Fixed RECAL connection and delays.
--  520730 - MCB yml update to remove IOIDRPTRAIN timing path.
--  532287 - Change default value of parameter CAL_CALIBRATION_MODE.
--  545576 - MEM_MDDR_ODS attribute update.
-------------------------------------------------------

----- CELL X_MCB -----

library IEEE;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

library simprim;
use simprim.VCOMPONENTS.all; 

library secureip; 
use secureip.all; 

use simprim.VPACKAGE.all;

  entity X_MCB is
    generic (
      TimingChecksOn : boolean := TRUE;
      InstancePath   : string  := "*";
      Xon            : boolean := TRUE;
      MsgOn          : boolean := FALSE;
      LOC            : string  := "UNPLACED";
      ARB_NUM_TIME_SLOTS : integer := 12;
      ARB_TIME_SLOT_0 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_1 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_10 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_11 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_2 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_3 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_4 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_5 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_6 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_7 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_8 : bit_vector := "111111111111111111";
      ARB_TIME_SLOT_9 : bit_vector := "111111111111111111";
      CAL_BA : bit_vector := X"0";
      CAL_BYPASS : string := "YES";
      CAL_CA : bit_vector := X"000";
      CAL_CALIBRATION_MODE : string := "NOCALIBRATION";
      CAL_CLK_DIV : integer := 1;
      CAL_DELAY : string := "QUARTER";
      CAL_RA : bit_vector := X"0000";
      MEM_ADDR_ORDER : string := "BANK_ROW_COLUMN";
      MEM_BA_SIZE : integer := 3;
      MEM_BURST_LEN : integer := 8;
      MEM_CAS_LATENCY : integer := 4;
      MEM_CA_SIZE : integer := 11;
      MEM_DDR1_2_ODS : string := "FULL";
      MEM_DDR2_3_HIGH_TEMP_SR : string := "NORMAL";
      MEM_DDR2_3_PA_SR : string := "FULL";
      MEM_DDR2_ADD_LATENCY : integer := 0;
      MEM_DDR2_DIFF_DQS_EN : string := "YES";
      MEM_DDR2_RTT : string := "50OHMS";
      MEM_DDR2_WRT_RECOVERY : integer := 4;
      MEM_DDR3_ADD_LATENCY : string := "OFF";
      MEM_DDR3_AUTO_SR : string := "ENABLED";
      MEM_DDR3_CAS_LATENCY : integer := 7;
      MEM_DDR3_CAS_WR_LATENCY : integer := 5;
      MEM_DDR3_DYN_WRT_ODT : string := "OFF";
      MEM_DDR3_ODS : string := "DIV7";
      MEM_DDR3_RTT : string := "DIV2";
      MEM_DDR3_WRT_RECOVERY : integer := 7;
      MEM_MDDR_ODS : string := "FULL";
      MEM_MOBILE_PA_SR : string := "FULL";
      MEM_MOBILE_TC_SR : integer := 0;
      MEM_RAS_VAL : integer := 0;
      MEM_RA_SIZE : integer := 13;
      MEM_RCD_VAL : integer := 1;
      MEM_REFI_VAL : integer := 0;
      MEM_RFC_VAL : integer := 0;
      MEM_RP_VAL : integer := 0;
      MEM_RTP_VAL : integer := 0;
      MEM_TYPE : string := "DDR3";
      MEM_WIDTH : integer := 4;
      MEM_WR_VAL : integer := 0;
      MEM_WTR_VAL : integer := 3;
      PORT_CONFIG : string := "B32_B32_B32_B32";
      tipd_DQI : VitalDelayArrayType01 (15 downto 0) := (others => (0 ps, 0 ps));
      tipd_DQSIOIN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_DQSIOIP : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_IOIDRPSDI : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0ARBEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0CMDBA : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0CMDBL : VitalDelayArrayType01 (5 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0CMDCA : VitalDelayArrayType01 (11 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0CMDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0CMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0CMDINSTR : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0CMDRA : VitalDelayArrayType01 (14 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0RDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0RDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0RWRMASK : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0WRCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P0WRDATA : VitalDelayArrayType01 (31 downto 0) := (others => (0 ps, 0 ps));
      tipd_P0WREN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1ARBEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1CMDBA : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1CMDBL : VitalDelayArrayType01 (5 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1CMDCA : VitalDelayArrayType01 (11 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1CMDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1CMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1CMDINSTR : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1CMDRA : VitalDelayArrayType01 (14 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1RDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1RDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1RWRMASK : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1WRCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P1WRDATA : VitalDelayArrayType01 (31 downto 0) := (others => (0 ps, 0 ps));
      tipd_P1WREN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P2ARBEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P2CLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P2CMDBA : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P2CMDBL : VitalDelayArrayType01 (5 downto 0) := (others => (0 ps, 0 ps));
      tipd_P2CMDCA : VitalDelayArrayType01 (11 downto 0) := (others => (0 ps, 0 ps));
      tipd_P2CMDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P2CMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P2CMDINSTR : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P2CMDRA : VitalDelayArrayType01 (14 downto 0) := (others => (0 ps, 0 ps));
      tipd_P2EN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P2WRDATA : VitalDelayArrayType01 (31 downto 0) := (others => (0 ps, 0 ps));
      tipd_P2WRMASK : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3ARBEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P3CLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P3CMDBA : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3CMDBL : VitalDelayArrayType01 (5 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3CMDCA : VitalDelayArrayType01 (11 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3CMDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P3CMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P3CMDINSTR : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3CMDRA : VitalDelayArrayType01 (14 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3EN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P3WRDATA : VitalDelayArrayType01 (31 downto 0) := (others => (0 ps, 0 ps));
      tipd_P3WRMASK : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4ARBEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P4CLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P4CMDBA : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4CMDBL : VitalDelayArrayType01 (5 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4CMDCA : VitalDelayArrayType01 (11 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4CMDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P4CMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P4CMDINSTR : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4CMDRA : VitalDelayArrayType01 (14 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4EN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P4WRDATA : VitalDelayArrayType01 (31 downto 0) := (others => (0 ps, 0 ps));
      tipd_P4WRMASK : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5ARBEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P5CLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P5CMDBA : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5CMDBL : VitalDelayArrayType01 (5 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5CMDCA : VitalDelayArrayType01 (11 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5CMDCLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P5CMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P5CMDINSTR : VitalDelayArrayType01 (2 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5CMDRA : VitalDelayArrayType01 (14 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5EN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_P5WRDATA : VitalDelayArrayType01 (31 downto 0) := (others => (0 ps, 0 ps));
      tipd_P5WRMASK : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_PLLCE : VitalDelayArrayType01 (1 downto 0) := (others => (0 ps, 0 ps));
      tipd_PLLCLK : VitalDelayArrayType01 (1 downto 0) := (others => (0 ps, 0 ps));
      tipd_PLLLOCK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_RECAL : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_SELFREFRESHENTER : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_SYSRST : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UDQSIOIN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UDQSIOIP : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIADD : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIADDR : VitalDelayArrayType01 (4 downto 0) := (others => (0 ps, 0 ps));
      tipd_UIBROADCAST : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UICLK : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UICMD : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UICMDEN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UICMDIN : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UICS : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIDONECAL : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIDQCOUNT : VitalDelayArrayType01 (3 downto 0) := (others => (0 ps, 0 ps));
      tipd_UIDQLOWERDEC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIDQLOWERINC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIDQUPPERDEC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIDQUPPERINC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIDRPUPDATE : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UILDQSDEC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UILDQSINC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIREAD : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UISDI : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIUDQSDEC : VitalDelayType01 :=  (0 ps, 0 ps);
      tipd_UIUDQSINC : VitalDelayType01 :=  (0 ps, 0 ps);
      tpd_P0CMDCLK_P0CMDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0CMDCLK_P0CMDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0RDCLK_P0RDCOUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P0RDCLK_P0RDDATA : VitalDelayArrayType01(31 downto 0) := (others => (0 ps, 0 ps));
      tpd_P0RDCLK_P0RDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0RDCLK_P0RDERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0RDCLK_P0RDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0RDCLK_P0RDOVERFLOW : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0WRCLK_P0WRCOUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P0WRCLK_P0WREMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0WRCLK_P0WRERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0WRCLK_P0WRFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P0WRCLK_P0WRUNDERRUN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1CMDCLK_P1CMDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1CMDCLK_P1CMDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1RDCLK_P1RDCOUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P1RDCLK_P1RDDATA : VitalDelayArrayType01(31 downto 0) := (others => (0 ps, 0 ps));
      tpd_P1RDCLK_P1RDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1RDCLK_P1RDERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1RDCLK_P1RDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1RDCLK_P1RDOVERFLOW : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1WRCLK_P1WRCOUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P1WRCLK_P1WREMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1WRCLK_P1WRERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1WRCLK_P1WRFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P1WRCLK_P1WRUNDERRUN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CLK_P2COUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P2CLK_P2EMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CLK_P2ERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CLK_P2FULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CLK_P2RDDATA : VitalDelayArrayType01(31 downto 0) := (others => (0 ps, 0 ps));
      tpd_P2CLK_P2RDOVERFLOW : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CLK_P2WRUNDERRUN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CMDCLK_P2CMDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P2CMDCLK_P2CMDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CLK_P3COUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P3CLK_P3EMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CLK_P3ERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CLK_P3FULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CLK_P3RDDATA : VitalDelayArrayType01(31 downto 0) := (others => (0 ps, 0 ps));
      tpd_P3CLK_P3RDOVERFLOW : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CLK_P3WRUNDERRUN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CMDCLK_P3CMDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P3CMDCLK_P3CMDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CLK_P4COUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P4CLK_P4EMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CLK_P4ERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CLK_P4FULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CLK_P4RDDATA : VitalDelayArrayType01(31 downto 0) := (others => (0 ps, 0 ps));
      tpd_P4CLK_P4RDOVERFLOW : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CLK_P4WRUNDERRUN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CMDCLK_P4CMDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P4CMDCLK_P4CMDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CLK_P5COUNT : VitalDelayArrayType01(6 downto 0) := (others => (0 ps, 0 ps));
      tpd_P5CLK_P5EMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CLK_P5ERROR : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CLK_P5FULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CLK_P5RDDATA : VitalDelayArrayType01(31 downto 0) := (others => (0 ps, 0 ps));
      tpd_P5CLK_P5RDOVERFLOW : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CLK_P5WRUNDERRUN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CMDCLK_P5CMDEMPTY : VitalDelayType01 := (0 ps, 0 ps);
      tpd_P5CMDCLK_P5CMDFULL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_PLLCLK_DQIOWEN0 : VitalDelayArrayType01(1 downto 0) := (others => (0 ps, 0 ps));
      tpd_PLLCLK_DQSIOWEN90N : VitalDelayArrayType01(1 downto 0) := (others => (0 ps, 0 ps));
      tpd_PLLCLK_DQSIOWEN90P : VitalDelayArrayType01(1 downto 0) := (others => (0 ps, 0 ps));
      tpd_PLLCLK_SELFREFRESHMODE : VitalDelayArrayType01(1 downto 0) := (others => (0 ps, 0 ps));
      tpd_UICLK_IOIDRPADD : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_IOIDRPADDR : VitalDelayArrayType01(4 downto 0) := (others => (0 ps, 0 ps));
      tpd_UICLK_IOIDRPBROADCAST : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_IOIDRPCLK : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_IOIDRPCS : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_IOIDRPSDO : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_IOIDRPUPDATE : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_UOCALSTART : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_UOCMDREADYIN : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_UODATA : VitalDelayArrayType01(7 downto 0) := (others => (0 ps, 0 ps));
      tpd_UICLK_UODATAVALID : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_UODONECAL : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_UOREFRSHFLAG : VitalDelayType01 := (0 ps, 0 ps);
      tpd_UICLK_UOSDO : VitalDelayType01 := (0 ps, 0 ps);
      thold_IOIDRPSDI_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_IOIDRPSDI_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P0ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P0ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P0CMDBA_P0CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P0CMDBA_P0CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P0CMDBL_P0CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P0CMDBL_P0CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P0CMDCA_P0CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P0CMDCA_P0CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P0CMDEN_P0CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P0CMDEN_P0CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P0CMDINSTR_P0CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P0CMDINSTR_P0CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P0CMDRA_P0CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P0CMDRA_P0CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P0RDEN_P0RDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P0RDEN_P0RDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P0RWRMASK_P0WRCLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P0RWRMASK_P0WRCLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P0WRDATA_P0WRCLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P0WRDATA_P0WRCLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P0WREN_P0WRCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P0WREN_P0WRCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P1ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P1ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P1CMDBA_P1CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P1CMDBA_P1CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P1CMDBL_P1CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P1CMDBL_P1CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P1CMDCA_P1CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P1CMDCA_P1CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P1CMDEN_P1CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P1CMDEN_P1CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P1CMDINSTR_P1CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P1CMDINSTR_P1CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P1CMDRA_P1CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P1CMDRA_P1CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P1RDEN_P1RDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P1RDEN_P1RDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P1RWRMASK_P1WRCLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P1RWRMASK_P1WRCLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P1WRDATA_P1WRCLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P1WRDATA_P1WRCLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P1WREN_P1WRCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P1WREN_P1WRCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P2ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P2ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P2CMDBA_P2CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P2CMDBA_P2CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P2CMDBL_P2CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P2CMDBL_P2CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P2CMDCA_P2CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P2CMDCA_P2CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P2CMDEN_P2CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P2CMDEN_P2CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P2CMDINSTR_P2CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P2CMDINSTR_P2CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P2CMDRA_P2CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P2CMDRA_P2CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P2EN_P2CLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P2EN_P2CLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P2WRDATA_P2CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P2WRDATA_P2CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P2WRMASK_P2CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P2WRMASK_P2CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P3ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P3ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P3CMDBA_P3CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P3CMDBA_P3CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P3CMDBL_P3CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P3CMDBL_P3CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P3CMDCA_P3CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P3CMDCA_P3CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P3CMDEN_P3CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P3CMDEN_P3CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P3CMDINSTR_P3CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P3CMDINSTR_P3CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P3CMDRA_P3CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P3CMDRA_P3CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P3EN_P3CLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P3EN_P3CLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P3WRDATA_P3CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P3WRDATA_P3CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P3WRMASK_P3CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P3WRMASK_P3CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P4ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P4ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P4CMDBA_P4CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P4CMDBA_P4CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P4CMDBL_P4CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P4CMDBL_P4CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P4CMDCA_P4CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P4CMDCA_P4CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P4CMDEN_P4CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P4CMDEN_P4CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P4CMDINSTR_P4CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P4CMDINSTR_P4CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P4CMDRA_P4CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P4CMDRA_P4CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P4EN_P4CLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P4EN_P4CLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P4WRDATA_P4CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P4WRDATA_P4CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P4WRMASK_P4CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P4WRMASK_P4CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P5ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P5ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_P5CMDBA_P5CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P5CMDBA_P5CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P5CMDBL_P5CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P5CMDBL_P5CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      thold_P5CMDCA_P5CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P5CMDCA_P5CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      thold_P5CMDEN_P5CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P5CMDEN_P5CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P5CMDINSTR_P5CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P5CMDINSTR_P5CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      thold_P5CMDRA_P5CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P5CMDRA_P5CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      thold_P5EN_P5CLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_P5EN_P5CLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_P5WRDATA_P5CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P5WRDATA_P5CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      thold_P5WRMASK_P5CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_P5WRMASK_P5CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_PLLCE_PLLCLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_PLLCE_PLLCLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_PLLLOCK_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_PLLLOCK_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_RECAL_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_RECAL_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_SELFREFRESHENTER_PLLCLK_negedge_negedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_SELFREFRESHENTER_PLLCLK_posedge_negedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      thold_UIADDR_UICLK_negedge_posedge : VitalDelayArrayType(4 downto 0) := (others => 0 ps);
      thold_UIADDR_UICLK_posedge_posedge : VitalDelayArrayType(4 downto 0) := (others => 0 ps);
      thold_UIADD_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIADD_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIBROADCAST_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIBROADCAST_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UICMDEN_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UICMDEN_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UICMDIN_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UICMDIN_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UICMD_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UICMD_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UICS_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UICS_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIDONECAL_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIDONECAL_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQCOUNT_UICLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_UIDQCOUNT_UICLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      thold_UIDQLOWERDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQLOWERDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQLOWERINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQLOWERINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQUPPERDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQUPPERDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQUPPERINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIDQUPPERINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIDRPUPDATE_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIDRPUPDATE_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UILDQSDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UILDQSDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UILDQSINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UILDQSINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIREAD_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIREAD_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UISDI_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UISDI_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIUDQSDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIUDQSDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      thold_UIUDQSINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      thold_UIUDQSINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_IOIDRPSDI_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_IOIDRPSDI_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P0ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P0ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P0CMDBA_P0CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P0CMDBA_P0CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P0CMDBL_P0CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P0CMDBL_P0CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P0CMDCA_P0CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P0CMDCA_P0CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P0CMDEN_P0CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P0CMDEN_P0CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P0CMDINSTR_P0CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P0CMDINSTR_P0CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P0CMDRA_P0CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P0CMDRA_P0CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P0RDEN_P0RDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P0RDEN_P0RDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P0RWRMASK_P0WRCLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P0RWRMASK_P0WRCLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P0WRDATA_P0WRCLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P0WRDATA_P0WRCLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P0WREN_P0WRCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P0WREN_P0WRCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P1ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P1ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P1CMDBA_P1CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P1CMDBA_P1CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P1CMDBL_P1CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P1CMDBL_P1CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P1CMDCA_P1CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P1CMDCA_P1CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P1CMDEN_P1CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P1CMDEN_P1CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P1CMDINSTR_P1CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P1CMDINSTR_P1CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P1CMDRA_P1CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P1CMDRA_P1CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P1RDEN_P1RDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P1RDEN_P1RDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P1RWRMASK_P1WRCLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P1RWRMASK_P1WRCLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P1WRDATA_P1WRCLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P1WRDATA_P1WRCLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P1WREN_P1WRCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P1WREN_P1WRCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P2ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P2ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P2CMDBA_P2CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P2CMDBA_P2CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P2CMDBL_P2CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P2CMDBL_P2CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P2CMDCA_P2CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P2CMDCA_P2CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P2CMDEN_P2CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P2CMDEN_P2CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P2CMDINSTR_P2CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P2CMDINSTR_P2CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P2CMDRA_P2CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P2CMDRA_P2CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P2EN_P2CLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P2EN_P2CLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P2WRDATA_P2CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P2WRDATA_P2CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P2WRMASK_P2CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P2WRMASK_P2CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P3ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P3ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P3CMDBA_P3CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P3CMDBA_P3CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P3CMDBL_P3CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P3CMDBL_P3CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P3CMDCA_P3CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P3CMDCA_P3CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P3CMDEN_P3CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P3CMDEN_P3CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P3CMDINSTR_P3CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P3CMDINSTR_P3CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P3CMDRA_P3CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P3CMDRA_P3CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P3EN_P3CLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P3EN_P3CLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P3WRDATA_P3CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P3WRDATA_P3CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P3WRMASK_P3CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P3WRMASK_P3CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P4ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P4ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P4CMDBA_P4CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P4CMDBA_P4CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P4CMDBL_P4CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P4CMDBL_P4CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P4CMDCA_P4CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P4CMDCA_P4CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P4CMDEN_P4CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P4CMDEN_P4CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P4CMDINSTR_P4CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P4CMDINSTR_P4CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P4CMDRA_P4CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P4CMDRA_P4CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P4EN_P4CLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P4EN_P4CLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P4WRDATA_P4CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P4WRDATA_P4CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P4WRMASK_P4CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P4WRMASK_P4CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P5ARBEN_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P5ARBEN_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_P5CMDBA_P5CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P5CMDBA_P5CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P5CMDBL_P5CMDCLK_negedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P5CMDBL_P5CMDCLK_posedge_posedge : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tsetup_P5CMDCA_P5CMDCLK_negedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P5CMDCA_P5CMDCLK_posedge_posedge : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tsetup_P5CMDEN_P5CMDCLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P5CMDEN_P5CMDCLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P5CMDINSTR_P5CMDCLK_negedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P5CMDINSTR_P5CMDCLK_posedge_posedge : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tsetup_P5CMDRA_P5CMDCLK_negedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P5CMDRA_P5CMDCLK_posedge_posedge : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tsetup_P5EN_P5CLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_P5EN_P5CLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_P5WRDATA_P5CLK_negedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P5WRDATA_P5CLK_posedge_posedge : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tsetup_P5WRMASK_P5CLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_P5WRMASK_P5CLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_PLLCE_PLLCLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_PLLCE_PLLCLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_PLLLOCK_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_PLLLOCK_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_RECAL_PLLCLK_negedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_RECAL_PLLCLK_posedge_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_SELFREFRESHENTER_PLLCLK_negedge_negedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_SELFREFRESHENTER_PLLCLK_posedge_negedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tsetup_UIADDR_UICLK_negedge_posedge : VitalDelayArrayType(4 downto 0) := (others => 0 ps);
      tsetup_UIADDR_UICLK_posedge_posedge : VitalDelayArrayType(4 downto 0) := (others => 0 ps);
      tsetup_UIADD_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIADD_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIBROADCAST_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIBROADCAST_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICMDEN_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICMDEN_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICMDIN_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICMDIN_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICMD_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICMD_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICS_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UICS_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDONECAL_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDONECAL_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQCOUNT_UICLK_negedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_UIDQCOUNT_UICLK_posedge_posedge : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tsetup_UIDQLOWERDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQLOWERDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQLOWERINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQLOWERINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQUPPERDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQUPPERDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQUPPERINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDQUPPERINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDRPUPDATE_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIDRPUPDATE_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UILDQSDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UILDQSDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UILDQSINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UILDQSINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIREAD_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIREAD_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UISDI_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UISDI_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIUDQSDEC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIUDQSDEC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIUDQSINC_UICLK_negedge_posedge : VitalDelayType := 0 ps;
      tsetup_UIUDQSINC_UICLK_posedge_posedge : VitalDelayType := 0 ps;
      tisd_IOIDRPSDI_UICLK : VitalDelayType := 0 ps;
      tisd_P0ARBEN_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_P0CMDBA_P0CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P0CMDBL_P0CMDCLK : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tisd_P0CMDCA_P0CMDCLK : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tisd_P0CMDEN_P0CMDCLK : VitalDelayType := 0 ps;
      tisd_P0CMDINSTR_P0CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P0CMDRA_P0CMDCLK : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tisd_P0RDEN_P0RDCLK : VitalDelayType := 0 ps;
      tisd_P0RWRMASK_P0WRCLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_P0WRDATA_P0WRCLK : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tisd_P0WREN_P0WRCLK : VitalDelayType := 0 ps;
      tisd_P1ARBEN_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_P1CMDBA_P1CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P1CMDBL_P1CMDCLK : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tisd_P1CMDCA_P1CMDCLK : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tisd_P1CMDEN_P1CMDCLK : VitalDelayType := 0 ps;
      tisd_P1CMDINSTR_P1CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P1CMDRA_P1CMDCLK : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tisd_P1RDEN_P1RDCLK : VitalDelayType := 0 ps;
      tisd_P1RWRMASK_P1WRCLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_P1WRDATA_P1WRCLK : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tisd_P1WREN_P1WRCLK : VitalDelayType := 0 ps;
      tisd_P2ARBEN_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_P2CMDBA_P2CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P2CMDBL_P2CMDCLK : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tisd_P2CMDCA_P2CMDCLK : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tisd_P2CMDEN_P2CMDCLK : VitalDelayType := 0 ps;
      tisd_P2CMDINSTR_P2CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P2CMDRA_P2CMDCLK : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tisd_P2EN_P2CLK : VitalDelayType := 0 ps;
      tisd_P2WRDATA_P2CLK : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tisd_P2WRMASK_P2CLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_P3ARBEN_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_P3CMDBA_P3CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P3CMDBL_P3CMDCLK : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tisd_P3CMDCA_P3CMDCLK : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tisd_P3CMDEN_P3CMDCLK : VitalDelayType := 0 ps;
      tisd_P3CMDINSTR_P3CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P3CMDRA_P3CMDCLK : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tisd_P3EN_P3CLK : VitalDelayType := 0 ps;
      tisd_P3WRDATA_P3CLK : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tisd_P3WRMASK_P3CLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_P4ARBEN_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_P4CMDBA_P4CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P4CMDBL_P4CMDCLK : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tisd_P4CMDCA_P4CMDCLK : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tisd_P4CMDEN_P4CMDCLK : VitalDelayType := 0 ps;
      tisd_P4CMDINSTR_P4CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P4CMDRA_P4CMDCLK : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tisd_P4EN_P4CLK : VitalDelayType := 0 ps;
      tisd_P4WRDATA_P4CLK : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tisd_P4WRMASK_P4CLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_P5ARBEN_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_P5CMDBA_P5CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P5CMDBL_P5CMDCLK : VitalDelayArrayType(5 downto 0) := (others => 0 ps);
      tisd_P5CMDCA_P5CMDCLK : VitalDelayArrayType(11 downto 0) := (others => 0 ps);
      tisd_P5CMDEN_P5CMDCLK : VitalDelayType := 0 ps;
      tisd_P5CMDINSTR_P5CMDCLK : VitalDelayArrayType(2 downto 0) := (others => 0 ps);
      tisd_P5CMDRA_P5CMDCLK : VitalDelayArrayType(14 downto 0) := (others => 0 ps);
      tisd_P5EN_P5CLK : VitalDelayType := 0 ps;
      tisd_P5WRDATA_P5CLK : VitalDelayArrayType(31 downto 0) := (others => 0 ps);
      tisd_P5WRMASK_P5CLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_PLLCE_PLLCLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_PLLLOCK_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_RECAL_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_SELFREFRESHENTER_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tisd_UIADDR_UICLK : VitalDelayArrayType(4 downto 0) := (others => 0 ps);
      tisd_UIADD_UICLK : VitalDelayType := 0 ps;
      tisd_UIBROADCAST_UICLK : VitalDelayType := 0 ps;
      tisd_UICMDEN_UICLK : VitalDelayType := 0 ps;
      tisd_UICMDIN_UICLK : VitalDelayType := 0 ps;
      tisd_UICMD_UICLK : VitalDelayType := 0 ps;
      tisd_UICS_UICLK : VitalDelayType := 0 ps;
      tisd_UIDONECAL_UICLK : VitalDelayType := 0 ps;
      tisd_UIDQCOUNT_UICLK : VitalDelayArrayType(3 downto 0) := (others => 0 ps);
      tisd_UIDQLOWERDEC_UICLK : VitalDelayType := 0 ps;
      tisd_UIDQLOWERINC_UICLK : VitalDelayType := 0 ps;
      tisd_UIDQUPPERDEC_UICLK : VitalDelayType := 0 ps;
      tisd_UIDQUPPERINC_UICLK : VitalDelayType := 0 ps;
      tisd_UIDRPUPDATE_UICLK : VitalDelayType := 0 ps;
      tisd_UILDQSDEC_UICLK : VitalDelayType := 0 ps;
      tisd_UILDQSINC_UICLK : VitalDelayType := 0 ps;
      tisd_UIREAD_UICLK : VitalDelayType := 0 ps;
      tisd_UISDI_UICLK : VitalDelayType := 0 ps;
      tisd_UIUDQSDEC_UICLK : VitalDelayType := 0 ps;
      tisd_UIUDQSINC_UICLK : VitalDelayType := 0 ps;
      ticd_P0CMDCLK : VitalDelayType := 0 ps;
      ticd_P0RDCLK : VitalDelayType := 0 ps;
      ticd_P0WRCLK : VitalDelayType := 0 ps;
      ticd_P1CMDCLK : VitalDelayType := 0 ps;
      ticd_P1RDCLK : VitalDelayType := 0 ps;
      ticd_P1WRCLK : VitalDelayType := 0 ps;
      ticd_P2CLK : VitalDelayType := 0 ps;
      ticd_P2CMDCLK : VitalDelayType := 0 ps;
      ticd_P3CLK : VitalDelayType := 0 ps;
      ticd_P3CMDCLK : VitalDelayType := 0 ps;
      ticd_P4CLK : VitalDelayType := 0 ps;
      ticd_P4CMDCLK : VitalDelayType := 0 ps;
      ticd_P5CLK : VitalDelayType := 0 ps;
      ticd_P5CMDCLK : VitalDelayType := 0 ps;
      ticd_PLLCLK : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      ticd_UICLK : VitalDelayType := 0 ps;
      tperiod_P0CMDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P0RDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P0WRCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P1CMDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P1RDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P1WRCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P2CLK_posedge : VitalDelayType := 0 ps;
      tperiod_P2CMDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P3CLK_posedge : VitalDelayType := 0 ps;
      tperiod_P3CMDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P4CLK_posedge : VitalDelayType := 0 ps;
      tperiod_P4CMDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_P5CLK_posedge : VitalDelayType := 0 ps;
      tperiod_P5CMDCLK_posedge : VitalDelayType := 0 ps;
      tperiod_PLLCLK_posedge : VitalDelayArrayType(1 downto 0) := (others => 0 ps);
      tperiod_SYSRST_posedge : VitalDelayType := 0 ps;
      tperiod_UICLK_posedge : VitalDelayType := 0 ps
    );

    port (
      ADDR                 : out std_logic_vector(14 downto 0);
      BA                   : out std_logic_vector(2 downto 0);
      CAS                  : out std_ulogic;
      CKE                  : out std_ulogic;
      DQIOWEN0             : out std_ulogic;
      DQON                 : out std_logic_vector(15 downto 0);
      DQOP                 : out std_logic_vector(15 downto 0);
      DQSIOWEN90N          : out std_ulogic;
      DQSIOWEN90P          : out std_ulogic;
      IOIDRPADD            : out std_ulogic;
      IOIDRPADDR           : out std_logic_vector(4 downto 0);
      IOIDRPBROADCAST      : out std_ulogic;
      IOIDRPCLK            : out std_ulogic;
      IOIDRPCS             : out std_ulogic;
      IOIDRPSDO            : out std_ulogic;
      IOIDRPTRAIN          : out std_ulogic;
      IOIDRPUPDATE         : out std_ulogic;
      LDMN                 : out std_ulogic;
      LDMP                 : out std_ulogic;
      ODT                  : out std_ulogic;
      P0CMDEMPTY           : out std_ulogic;
      P0CMDFULL            : out std_ulogic;
      P0RDCOUNT            : out std_logic_vector(6 downto 0);
      P0RDDATA             : out std_logic_vector(31 downto 0);
      P0RDEMPTY            : out std_ulogic;
      P0RDERROR            : out std_ulogic;
      P0RDFULL             : out std_ulogic;
      P0RDOVERFLOW         : out std_ulogic;
      P0WRCOUNT            : out std_logic_vector(6 downto 0);
      P0WREMPTY            : out std_ulogic;
      P0WRERROR            : out std_ulogic;
      P0WRFULL             : out std_ulogic;
      P0WRUNDERRUN         : out std_ulogic;
      P1CMDEMPTY           : out std_ulogic;
      P1CMDFULL            : out std_ulogic;
      P1RDCOUNT            : out std_logic_vector(6 downto 0);
      P1RDDATA             : out std_logic_vector(31 downto 0);
      P1RDEMPTY            : out std_ulogic;
      P1RDERROR            : out std_ulogic;
      P1RDFULL             : out std_ulogic;
      P1RDOVERFLOW         : out std_ulogic;
      P1WRCOUNT            : out std_logic_vector(6 downto 0);
      P1WREMPTY            : out std_ulogic;
      P1WRERROR            : out std_ulogic;
      P1WRFULL             : out std_ulogic;
      P1WRUNDERRUN         : out std_ulogic;
      P2CMDEMPTY           : out std_ulogic;
      P2CMDFULL            : out std_ulogic;
      P2COUNT              : out std_logic_vector(6 downto 0);
      P2EMPTY              : out std_ulogic;
      P2ERROR              : out std_ulogic;
      P2FULL               : out std_ulogic;
      P2RDDATA             : out std_logic_vector(31 downto 0);
      P2RDOVERFLOW         : out std_ulogic;
      P2WRUNDERRUN         : out std_ulogic;
      P3CMDEMPTY           : out std_ulogic;
      P3CMDFULL            : out std_ulogic;
      P3COUNT              : out std_logic_vector(6 downto 0);
      P3EMPTY              : out std_ulogic;
      P3ERROR              : out std_ulogic;
      P3FULL               : out std_ulogic;
      P3RDDATA             : out std_logic_vector(31 downto 0);
      P3RDOVERFLOW         : out std_ulogic;
      P3WRUNDERRUN         : out std_ulogic;
      P4CMDEMPTY           : out std_ulogic;
      P4CMDFULL            : out std_ulogic;
      P4COUNT              : out std_logic_vector(6 downto 0);
      P4EMPTY              : out std_ulogic;
      P4ERROR              : out std_ulogic;
      P4FULL               : out std_ulogic;
      P4RDDATA             : out std_logic_vector(31 downto 0);
      P4RDOVERFLOW         : out std_ulogic;
      P4WRUNDERRUN         : out std_ulogic;
      P5CMDEMPTY           : out std_ulogic;
      P5CMDFULL            : out std_ulogic;
      P5COUNT              : out std_logic_vector(6 downto 0);
      P5EMPTY              : out std_ulogic;
      P5ERROR              : out std_ulogic;
      P5FULL               : out std_ulogic;
      P5RDDATA             : out std_logic_vector(31 downto 0);
      P5RDOVERFLOW         : out std_ulogic;
      P5WRUNDERRUN         : out std_ulogic;
      RAS                  : out std_ulogic;
      RST                  : out std_ulogic;
      SELFREFRESHMODE      : out std_ulogic;
      STATUS               : out std_logic_vector(31 downto 0);
      UDMN                 : out std_ulogic;
      UDMP                 : out std_ulogic;
      UOCALSTART           : out std_ulogic;
      UOCMDREADYIN         : out std_ulogic;
      UODATA               : out std_logic_vector(7 downto 0);
      UODATAVALID          : out std_ulogic;
      UODONECAL            : out std_ulogic;
      UOREFRSHFLAG         : out std_ulogic;
      UOSDO                : out std_ulogic;
      WE                   : out std_ulogic;
      DQI                  : in std_logic_vector(15 downto 0);
      DQSIOIN              : in std_ulogic;
      DQSIOIP              : in std_ulogic;
      IOIDRPSDI            : in std_ulogic;
      P0ARBEN              : in std_ulogic;
      P0CMDBA              : in std_logic_vector(2 downto 0);
      P0CMDBL              : in std_logic_vector(5 downto 0);
      P0CMDCA              : in std_logic_vector(11 downto 0);
      P0CMDCLK             : in std_ulogic;
      P0CMDEN              : in std_ulogic;
      P0CMDINSTR           : in std_logic_vector(2 downto 0);
      P0CMDRA              : in std_logic_vector(14 downto 0);
      P0RDCLK              : in std_ulogic;
      P0RDEN               : in std_ulogic;
      P0RWRMASK            : in std_logic_vector(3 downto 0);
      P0WRCLK              : in std_ulogic;
      P0WRDATA             : in std_logic_vector(31 downto 0);
      P0WREN               : in std_ulogic;
      P1ARBEN              : in std_ulogic;
      P1CMDBA              : in std_logic_vector(2 downto 0);
      P1CMDBL              : in std_logic_vector(5 downto 0);
      P1CMDCA              : in std_logic_vector(11 downto 0);
      P1CMDCLK             : in std_ulogic;
      P1CMDEN              : in std_ulogic;
      P1CMDINSTR           : in std_logic_vector(2 downto 0);
      P1CMDRA              : in std_logic_vector(14 downto 0);
      P1RDCLK              : in std_ulogic;
      P1RDEN               : in std_ulogic;
      P1RWRMASK            : in std_logic_vector(3 downto 0);
      P1WRCLK              : in std_ulogic;
      P1WRDATA             : in std_logic_vector(31 downto 0);
      P1WREN               : in std_ulogic;
      P2ARBEN              : in std_ulogic;
      P2CLK                : in std_ulogic;
      P2CMDBA              : in std_logic_vector(2 downto 0);
      P2CMDBL              : in std_logic_vector(5 downto 0);
      P2CMDCA              : in std_logic_vector(11 downto 0);
      P2CMDCLK             : in std_ulogic;
      P2CMDEN              : in std_ulogic;
      P2CMDINSTR           : in std_logic_vector(2 downto 0);
      P2CMDRA              : in std_logic_vector(14 downto 0);
      P2EN                 : in std_ulogic;
      P2WRDATA             : in std_logic_vector(31 downto 0);
      P2WRMASK             : in std_logic_vector(3 downto 0);
      P3ARBEN              : in std_ulogic;
      P3CLK                : in std_ulogic;
      P3CMDBA              : in std_logic_vector(2 downto 0);
      P3CMDBL              : in std_logic_vector(5 downto 0);
      P3CMDCA              : in std_logic_vector(11 downto 0);
      P3CMDCLK             : in std_ulogic;
      P3CMDEN              : in std_ulogic;
      P3CMDINSTR           : in std_logic_vector(2 downto 0);
      P3CMDRA              : in std_logic_vector(14 downto 0);
      P3EN                 : in std_ulogic;
      P3WRDATA             : in std_logic_vector(31 downto 0);
      P3WRMASK             : in std_logic_vector(3 downto 0);
      P4ARBEN              : in std_ulogic;
      P4CLK                : in std_ulogic;
      P4CMDBA              : in std_logic_vector(2 downto 0);
      P4CMDBL              : in std_logic_vector(5 downto 0);
      P4CMDCA              : in std_logic_vector(11 downto 0);
      P4CMDCLK             : in std_ulogic;
      P4CMDEN              : in std_ulogic;
      P4CMDINSTR           : in std_logic_vector(2 downto 0);
      P4CMDRA              : in std_logic_vector(14 downto 0);
      P4EN                 : in std_ulogic;
      P4WRDATA             : in std_logic_vector(31 downto 0);
      P4WRMASK             : in std_logic_vector(3 downto 0);
      P5ARBEN              : in std_ulogic;
      P5CLK                : in std_ulogic;
      P5CMDBA              : in std_logic_vector(2 downto 0);
      P5CMDBL              : in std_logic_vector(5 downto 0);
      P5CMDCA              : in std_logic_vector(11 downto 0);
      P5CMDCLK             : in std_ulogic;
      P5CMDEN              : in std_ulogic;
      P5CMDINSTR           : in std_logic_vector(2 downto 0);
      P5CMDRA              : in std_logic_vector(14 downto 0);
      P5EN                 : in std_ulogic;
      P5WRDATA             : in std_logic_vector(31 downto 0);
      P5WRMASK             : in std_logic_vector(3 downto 0);
      PLLCE                : in std_logic_vector(1 downto 0);
      PLLCLK               : in std_logic_vector(1 downto 0);
      PLLLOCK              : in std_ulogic;
      RECAL                : in std_ulogic;
      SELFREFRESHENTER     : in std_ulogic;
      SYSRST               : in std_ulogic;
      UDQSIOIN             : in std_ulogic;
      UDQSIOIP             : in std_ulogic;
      UIADD                : in std_ulogic;
      UIADDR               : in std_logic_vector(4 downto 0);
      UIBROADCAST          : in std_ulogic;
      UICLK                : in std_ulogic;
      UICMD                : in std_ulogic;
      UICMDEN              : in std_ulogic;
      UICMDIN              : in std_ulogic;
      UICS                 : in std_ulogic;
      UIDONECAL            : in std_ulogic;
      UIDQCOUNT            : in std_logic_vector(3 downto 0);
      UIDQLOWERDEC         : in std_ulogic;
      UIDQLOWERINC         : in std_ulogic;
      UIDQUPPERDEC         : in std_ulogic;
      UIDQUPPERINC         : in std_ulogic;
      UIDRPUPDATE          : in std_ulogic;
      UILDQSDEC            : in std_ulogic;
      UILDQSINC            : in std_ulogic;
      UIREAD               : in std_ulogic;
      UISDI                : in std_ulogic;
      UIUDQSDEC            : in std_ulogic;
      UIUDQSINC            : in std_ulogic      
    );
    attribute VITAL_LEVEL0 of X_MCB :     entity is true;
  end X_MCB;

  architecture X_MCB_V of X_MCB is
    TYPE VitalTimingDataArrayType IS ARRAY (NATURAL RANGE <>) OF VitalTimingDataType;
    component MCB_WRAP
      generic (
        ARB_NUM_TIME_SLOTS : integer;
        ARB_TIME_SLOT_0 : string;
        ARB_TIME_SLOT_1 : string;
        ARB_TIME_SLOT_10 : string;
        ARB_TIME_SLOT_11 : string;
        ARB_TIME_SLOT_2 : string;
        ARB_TIME_SLOT_3 : string;
        ARB_TIME_SLOT_4 : string;
        ARB_TIME_SLOT_5 : string;
        ARB_TIME_SLOT_6 : string;
        ARB_TIME_SLOT_7 : string;
        ARB_TIME_SLOT_8 : string;
        ARB_TIME_SLOT_9 : string;
        CAL_BA : string;
        CAL_BYPASS : string;
        CAL_CA : string;
        CAL_CALIBRATION_MODE : string;
        CAL_CLK_DIV : integer;
        CAL_DELAY : string;
        CAL_RA : string;
        MEM_ADDR_ORDER : string;
        MEM_BA_SIZE : integer;
        MEM_BURST_LEN : integer;
        MEM_CAS_LATENCY : integer;
        MEM_CA_SIZE : integer;
        MEM_DDR1_2_ODS : string;
        MEM_DDR2_3_HIGH_TEMP_SR : string;
        MEM_DDR2_3_PA_SR : string;
        MEM_DDR2_ADD_LATENCY : integer;
        MEM_DDR2_DIFF_DQS_EN : string;
        MEM_DDR2_RTT : string;
        MEM_DDR2_WRT_RECOVERY : integer;
        MEM_DDR3_ADD_LATENCY : string;
        MEM_DDR3_AUTO_SR : string;
        MEM_DDR3_CAS_LATENCY : integer;
        MEM_DDR3_CAS_WR_LATENCY : integer;
        MEM_DDR3_DYN_WRT_ODT : string;
        MEM_DDR3_ODS : string;
        MEM_DDR3_RTT : string;
        MEM_DDR3_WRT_RECOVERY : integer;
        MEM_MDDR_ODS : string;
        MEM_MOBILE_PA_SR : string;
        MEM_MOBILE_TC_SR : integer;
        MEM_RAS_VAL : integer;
        MEM_RA_SIZE : integer;
        MEM_RCD_VAL : integer;
        MEM_REFI_VAL : integer;
        MEM_RFC_VAL : integer;
        MEM_RP_VAL : integer;
        MEM_RTP_VAL : integer;
        MEM_TYPE : string;
        MEM_WIDTH : integer;
        MEM_WR_VAL : integer;
        MEM_WTR_VAL : integer;
        PORT_CONFIG : string        
      );
      
      port (
        ADDR                 : out std_logic_vector(14 downto 0);
        BA                   : out std_logic_vector(2 downto 0);
        CAS                  : out std_ulogic;
        CKE                  : out std_ulogic;
        DQIOWEN0             : out std_ulogic;
        DQON                 : out std_logic_vector(15 downto 0);
        DQOP                 : out std_logic_vector(15 downto 0);
        DQSIOWEN90N          : out std_ulogic;
        DQSIOWEN90P          : out std_ulogic;
        IOIDRPADD            : out std_ulogic;
        IOIDRPADDR           : out std_logic_vector(4 downto 0);
        IOIDRPBROADCAST      : out std_ulogic;
        IOIDRPCLK            : out std_ulogic;
        IOIDRPCS             : out std_ulogic;
        IOIDRPSDO            : out std_ulogic;
        IOIDRPTRAIN          : out std_ulogic;
        IOIDRPUPDATE         : out std_ulogic;
        LDMN                 : out std_ulogic;
        LDMP                 : out std_ulogic;
        ODT                  : out std_ulogic;
        P0CMDEMPTY           : out std_ulogic;
        P0CMDFULL            : out std_ulogic;
        P0RDCOUNT            : out std_logic_vector(6 downto 0);
        P0RDDATA             : out std_logic_vector(31 downto 0);
        P0RDEMPTY            : out std_ulogic;
        P0RDERROR            : out std_ulogic;
        P0RDFULL             : out std_ulogic;
        P0RDOVERFLOW         : out std_ulogic;
        P0WRCOUNT            : out std_logic_vector(6 downto 0);
        P0WREMPTY            : out std_ulogic;
        P0WRERROR            : out std_ulogic;
        P0WRFULL             : out std_ulogic;
        P0WRUNDERRUN         : out std_ulogic;
        P1CMDEMPTY           : out std_ulogic;
        P1CMDFULL            : out std_ulogic;
        P1RDCOUNT            : out std_logic_vector(6 downto 0);
        P1RDDATA             : out std_logic_vector(31 downto 0);
        P1RDEMPTY            : out std_ulogic;
        P1RDERROR            : out std_ulogic;
        P1RDFULL             : out std_ulogic;
        P1RDOVERFLOW         : out std_ulogic;
        P1WRCOUNT            : out std_logic_vector(6 downto 0);
        P1WREMPTY            : out std_ulogic;
        P1WRERROR            : out std_ulogic;
        P1WRFULL             : out std_ulogic;
        P1WRUNDERRUN         : out std_ulogic;
        P2CMDEMPTY           : out std_ulogic;
        P2CMDFULL            : out std_ulogic;
        P2COUNT              : out std_logic_vector(6 downto 0);
        P2EMPTY              : out std_ulogic;
        P2ERROR              : out std_ulogic;
        P2FULL               : out std_ulogic;
        P2RDDATA             : out std_logic_vector(31 downto 0);
        P2RDOVERFLOW         : out std_ulogic;
        P2WRUNDERRUN         : out std_ulogic;
        P3CMDEMPTY           : out std_ulogic;
        P3CMDFULL            : out std_ulogic;
        P3COUNT              : out std_logic_vector(6 downto 0);
        P3EMPTY              : out std_ulogic;
        P3ERROR              : out std_ulogic;
        P3FULL               : out std_ulogic;
        P3RDDATA             : out std_logic_vector(31 downto 0);
        P3RDOVERFLOW         : out std_ulogic;
        P3WRUNDERRUN         : out std_ulogic;
        P4CMDEMPTY           : out std_ulogic;
        P4CMDFULL            : out std_ulogic;
        P4COUNT              : out std_logic_vector(6 downto 0);
        P4EMPTY              : out std_ulogic;
        P4ERROR              : out std_ulogic;
        P4FULL               : out std_ulogic;
        P4RDDATA             : out std_logic_vector(31 downto 0);
        P4RDOVERFLOW         : out std_ulogic;
        P4WRUNDERRUN         : out std_ulogic;
        P5CMDEMPTY           : out std_ulogic;
        P5CMDFULL            : out std_ulogic;
        P5COUNT              : out std_logic_vector(6 downto 0);
        P5EMPTY              : out std_ulogic;
        P5ERROR              : out std_ulogic;
        P5FULL               : out std_ulogic;
        P5RDDATA             : out std_logic_vector(31 downto 0);
        P5RDOVERFLOW         : out std_ulogic;
        P5WRUNDERRUN         : out std_ulogic;
        RAS                  : out std_ulogic;
        RST                  : out std_ulogic;
        SELFREFRESHMODE      : out std_ulogic;
        STATUS               : out std_logic_vector(31 downto 0);
        UDMN                 : out std_ulogic;
        UDMP                 : out std_ulogic;
        UOCALSTART           : out std_ulogic;
        UOCMDREADYIN         : out std_ulogic;
        UODATA               : out std_logic_vector(7 downto 0);
        UODATAVALID          : out std_ulogic;
        UODONECAL            : out std_ulogic;
        UOREFRSHFLAG         : out std_ulogic;
        UOSDO                : out std_ulogic;
        WE                   : out std_ulogic;
        DQI                  : in std_logic_vector(15 downto 0);
        DQSIOIN              : in std_ulogic;
        DQSIOIP              : in std_ulogic;
        IOIDRPSDI            : in std_ulogic;
        P0ARBEN              : in std_ulogic;
        P0CMDBA              : in std_logic_vector(2 downto 0);
        P0CMDBL              : in std_logic_vector(5 downto 0);
        P0CMDCA              : in std_logic_vector(11 downto 0);
        P0CMDCLK             : in std_ulogic;
        P0CMDEN              : in std_ulogic;
        P0CMDINSTR           : in std_logic_vector(2 downto 0);
        P0CMDRA              : in std_logic_vector(14 downto 0);
        P0RDCLK              : in std_ulogic;
        P0RDEN               : in std_ulogic;
        P0RWRMASK            : in std_logic_vector(3 downto 0);
        P0WRCLK              : in std_ulogic;
        P0WRDATA             : in std_logic_vector(31 downto 0);
        P0WREN               : in std_ulogic;
        P1ARBEN              : in std_ulogic;
        P1CMDBA              : in std_logic_vector(2 downto 0);
        P1CMDBL              : in std_logic_vector(5 downto 0);
        P1CMDCA              : in std_logic_vector(11 downto 0);
        P1CMDCLK             : in std_ulogic;
        P1CMDEN              : in std_ulogic;
        P1CMDINSTR           : in std_logic_vector(2 downto 0);
        P1CMDRA              : in std_logic_vector(14 downto 0);
        P1RDCLK              : in std_ulogic;
        P1RDEN               : in std_ulogic;
        P1RWRMASK            : in std_logic_vector(3 downto 0);
        P1WRCLK              : in std_ulogic;
        P1WRDATA             : in std_logic_vector(31 downto 0);
        P1WREN               : in std_ulogic;
        P2ARBEN              : in std_ulogic;
        P2CLK                : in std_ulogic;
        P2CMDBA              : in std_logic_vector(2 downto 0);
        P2CMDBL              : in std_logic_vector(5 downto 0);
        P2CMDCA              : in std_logic_vector(11 downto 0);
        P2CMDCLK             : in std_ulogic;
        P2CMDEN              : in std_ulogic;
        P2CMDINSTR           : in std_logic_vector(2 downto 0);
        P2CMDRA              : in std_logic_vector(14 downto 0);
        P2EN                 : in std_ulogic;
        P2WRDATA             : in std_logic_vector(31 downto 0);
        P2WRMASK             : in std_logic_vector(3 downto 0);
        P3ARBEN              : in std_ulogic;
        P3CLK                : in std_ulogic;
        P3CMDBA              : in std_logic_vector(2 downto 0);
        P3CMDBL              : in std_logic_vector(5 downto 0);
        P3CMDCA              : in std_logic_vector(11 downto 0);
        P3CMDCLK             : in std_ulogic;
        P3CMDEN              : in std_ulogic;
        P3CMDINSTR           : in std_logic_vector(2 downto 0);
        P3CMDRA              : in std_logic_vector(14 downto 0);
        P3EN                 : in std_ulogic;
        P3WRDATA             : in std_logic_vector(31 downto 0);
        P3WRMASK             : in std_logic_vector(3 downto 0);
        P4ARBEN              : in std_ulogic;
        P4CLK                : in std_ulogic;
        P4CMDBA              : in std_logic_vector(2 downto 0);
        P4CMDBL              : in std_logic_vector(5 downto 0);
        P4CMDCA              : in std_logic_vector(11 downto 0);
        P4CMDCLK             : in std_ulogic;
        P4CMDEN              : in std_ulogic;
        P4CMDINSTR           : in std_logic_vector(2 downto 0);
        P4CMDRA              : in std_logic_vector(14 downto 0);
        P4EN                 : in std_ulogic;
        P4WRDATA             : in std_logic_vector(31 downto 0);
        P4WRMASK             : in std_logic_vector(3 downto 0);
        P5ARBEN              : in std_ulogic;
        P5CLK                : in std_ulogic;
        P5CMDBA              : in std_logic_vector(2 downto 0);
        P5CMDBL              : in std_logic_vector(5 downto 0);
        P5CMDCA              : in std_logic_vector(11 downto 0);
        P5CMDCLK             : in std_ulogic;
        P5CMDEN              : in std_ulogic;
        P5CMDINSTR           : in std_logic_vector(2 downto 0);
        P5CMDRA              : in std_logic_vector(14 downto 0);
        P5EN                 : in std_ulogic;
        P5WRDATA             : in std_logic_vector(31 downto 0);
        P5WRMASK             : in std_logic_vector(3 downto 0);
        PLLCE                : in std_logic_vector(1 downto 0);
        PLLCLK               : in std_logic_vector(1 downto 0);
        PLLLOCK              : in std_ulogic;
        RECAL                : in std_ulogic;
        SELFREFRESHENTER     : in std_ulogic;
        SYSRST               : in std_ulogic;
        UDQSIOIN             : in std_ulogic;
        UDQSIOIP             : in std_ulogic;
        UIADD                : in std_ulogic;
        UIADDR               : in std_logic_vector(4 downto 0);
        UIBROADCAST          : in std_ulogic;
        UICLK                : in std_ulogic;
        UICMD                : in std_ulogic;
        UICMDEN              : in std_ulogic;
        UICMDIN              : in std_ulogic;
        UICS                 : in std_ulogic;
        UIDONECAL            : in std_ulogic;
        UIDQCOUNT            : in std_logic_vector(3 downto 0);
        UIDQLOWERDEC         : in std_ulogic;
        UIDQLOWERINC         : in std_ulogic;
        UIDQUPPERDEC         : in std_ulogic;
        UIDQUPPERINC         : in std_ulogic;
        UIDRPUPDATE          : in std_ulogic;
        UILDQSDEC            : in std_ulogic;
        UILDQSINC            : in std_ulogic;
        UIREAD               : in std_ulogic;
        UISDI                : in std_ulogic;
        UIUDQSDEC            : in std_ulogic;
        UIUDQSINC            : in std_ulogic;        
        GSR                  : in std_ulogic
      );
    end component;
    
    constant IN_DELAY : time := 0 ps;
    constant OUT_DELAY : time := 100 ps;
    constant INCLK_DELAY : time := 0 ps;
    constant OUTCLK_DELAY : time := 100 ps;

    function boolean_to_string(bool: boolean)
    return string is
    begin
      if bool then
        return "TRUE";
      else
        return "FALSE";
      end if;
    end boolean_to_string;

    function getstrlength (
           in_vec : std_logic_vector)
    return integer is
     variable string_length : integer;
    begin
     if ((in_vec'length mod 4) = 0) then
      string_length := in_vec'length/4;
    elsif ((in_vec'length mod 4) > 0) then
      string_length := in_vec'length/4 + 1;
    end if;
    return string_length;
    end getstrlength;

    -- Convert bit_vector to std_logic_vector
    constant ARB_TIME_SLOT_0_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_0)(17 downto 0);
    constant ARB_TIME_SLOT_10_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_10)(17 downto 0);
    constant ARB_TIME_SLOT_11_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_11)(17 downto 0);
    constant ARB_TIME_SLOT_1_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_1)(17 downto 0);
    constant ARB_TIME_SLOT_2_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_2)(17 downto 0);
    constant ARB_TIME_SLOT_3_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_3)(17 downto 0);
    constant ARB_TIME_SLOT_4_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_4)(17 downto 0);
    constant ARB_TIME_SLOT_5_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_5)(17 downto 0);
    constant ARB_TIME_SLOT_6_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_6)(17 downto 0);
    constant ARB_TIME_SLOT_7_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_7)(17 downto 0);
    constant ARB_TIME_SLOT_8_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_8)(17 downto 0);
    constant ARB_TIME_SLOT_9_BINARY : std_logic_vector(17 downto 0) := To_StdLogicVector(ARB_TIME_SLOT_9)(17 downto 0);
    constant CAL_BA_BINARY : std_logic_vector(2 downto 0) := To_StdLogicVector(CAL_BA)(2 downto 0);
    constant CAL_CA_BINARY : std_logic_vector(11 downto 0) := To_StdLogicVector(CAL_CA)(11 downto 0);
    constant CAL_RA_BINARY : std_logic_vector(14 downto 0) := To_StdLogicVector(CAL_RA)(14 downto 0);

    -- Get String Length
    constant CAL_BA_STRLEN : integer := getstrlength(CAL_BA_BINARY);
    constant CAL_CA_STRLEN : integer := getstrlength(CAL_CA_BINARY);
    constant CAL_RA_STRLEN : integer := getstrlength(CAL_RA_BINARY);
    
    -- Convert std_logic_vector to string
    constant ARB_TIME_SLOT_0_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_0_BINARY);
    constant ARB_TIME_SLOT_10_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_10_BINARY);
    constant ARB_TIME_SLOT_11_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_11_BINARY);
    constant ARB_TIME_SLOT_1_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_1_BINARY);
    constant ARB_TIME_SLOT_2_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_2_BINARY);
    constant ARB_TIME_SLOT_3_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_3_BINARY);
    constant ARB_TIME_SLOT_4_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_4_BINARY);
    constant ARB_TIME_SLOT_5_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_5_BINARY);
    constant ARB_TIME_SLOT_6_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_6_BINARY);
    constant ARB_TIME_SLOT_7_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_7_BINARY);
    constant ARB_TIME_SLOT_8_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_8_BINARY);
    constant ARB_TIME_SLOT_9_STRING : string := SLV_TO_STR(ARB_TIME_SLOT_9_BINARY);
    constant CAL_BA_STRING : string := SLV_TO_HEX(CAL_BA_BINARY, CAL_BA_STRLEN);
    constant CAL_CA_STRING : string := SLV_TO_HEX(CAL_CA_BINARY, CAL_CA_STRLEN);
    constant CAL_RA_STRING : string := SLV_TO_HEX(CAL_RA_BINARY, CAL_RA_STRLEN);
    
    signal ARB_NUM_TIME_SLOTS_BINARY : std_ulogic;
    signal CAL_BYPASS_BINARY : std_ulogic;
    signal CAL_CALIBRATION_MODE_BINARY : std_ulogic;
    signal CAL_CLK_DIV_BINARY : std_logic_vector(2 downto 0);
    signal CAL_DELAY_BINARY : std_logic_vector(1 downto 0);
    signal MEM_ADDR_ORDER_BINARY : std_ulogic;
    signal MEM_BA_SIZE_BINARY : std_ulogic;
    signal MEM_BURST_LEN_BINARY : std_logic_vector(2 downto 0);
    signal MEM_CAS_LATENCY_BINARY : std_logic_vector(2 downto 0);
    signal MEM_CA_SIZE_BINARY : std_logic_vector(1 downto 0);
    signal MEM_DDR1_2_ODS_BINARY : std_ulogic;
    signal MEM_DDR2_3_HIGH_TEMP_SR_BINARY : std_ulogic;
    signal MEM_DDR2_3_PA_SR_BINARY : std_logic_vector(2 downto 0);
    signal MEM_DDR2_ADD_LATENCY_BINARY : std_logic_vector(2 downto 0);
    signal MEM_DDR2_DIFF_DQS_EN_BINARY : std_ulogic;
    signal MEM_DDR2_RTT_BINARY : std_logic_vector(1 downto 0);
    signal MEM_DDR2_WRT_RECOVERY_BINARY : std_logic_vector(2 downto 0);
    signal MEM_DDR3_ADD_LATENCY_BINARY : std_logic_vector(1 downto 0);
    signal MEM_DDR3_AUTO_SR_BINARY : std_ulogic;
    signal MEM_DDR3_CAS_LATENCY_BINARY : std_logic_vector(3 downto 0);
    signal MEM_DDR3_CAS_WR_LATENCY_BINARY : std_logic_vector(2 downto 0);
    signal MEM_DDR3_DYN_WRT_ODT_BINARY : std_logic_vector(1 downto 0);
    signal MEM_DDR3_ODS_BINARY : std_logic_vector(1 downto 0);
    signal MEM_DDR3_RTT_BINARY : std_logic_vector(2 downto 0);
    signal MEM_DDR3_WRT_RECOVERY_BINARY : std_logic_vector(2 downto 0);
    signal MEM_MDDR_ODS_BINARY : std_logic_vector(2 downto 0);
    signal MEM_MOBILE_PA_SR_BINARY : std_logic_vector(2 downto 0);
    signal MEM_MOBILE_TC_SR_BINARY : std_logic_vector(1 downto 0);
    signal MEM_RAS_VAL_BINARY : std_logic_vector(4 downto 0);
    signal MEM_RA_SIZE_BINARY : std_logic_vector(1 downto 0);
    signal MEM_RCD_VAL_BINARY : std_logic_vector(2 downto 0);
    signal MEM_REFI_VAL_BINARY : std_logic_vector(11 downto 0);
    signal MEM_RFC_VAL_BINARY : std_logic_vector(7 downto 0);
    signal MEM_RP_VAL_BINARY : std_logic_vector(3 downto 0);
    signal MEM_RTP_VAL_BINARY : std_logic_vector(2 downto 0);
    signal MEM_TYPE_BINARY : std_logic_vector(2 downto 0);
    signal MEM_WIDTH_BINARY : std_logic_vector(1 downto 0);
    signal MEM_WR_VAL_BINARY : std_logic_vector(2 downto 0);
    signal MEM_WTR_VAL_BINARY : std_logic_vector(2 downto 0);
    signal PORT_CONFIG_BINARY : std_logic_vector(2 downto 0);
    
    signal ADDR_out : std_logic_vector(14 downto 0);
    signal BA_out : std_logic_vector(2 downto 0);
    signal CAS_out : std_ulogic;
    signal CKE_out : std_ulogic;
    signal DQIOWEN0_out : std_ulogic;
    signal DQON_out : std_logic_vector(15 downto 0);
    signal DQOP_out : std_logic_vector(15 downto 0);
    signal DQSIOWEN90N_out : std_ulogic;
    signal DQSIOWEN90P_out : std_ulogic;
    signal IOIDRPADDR_out : std_logic_vector(4 downto 0);
    signal IOIDRPADD_out : std_ulogic;
    signal IOIDRPBROADCAST_out : std_ulogic;
    signal IOIDRPCLK_out : std_ulogic;
    signal IOIDRPCS_out : std_ulogic;
    signal IOIDRPSDO_out : std_ulogic;
    signal IOIDRPTRAIN_out : std_ulogic;
    signal IOIDRPUPDATE_out : std_ulogic;
    signal LDMN_out : std_ulogic;
    signal LDMP_out : std_ulogic;
    signal ODT_out : std_ulogic;
    signal P0CMDEMPTY_out : std_ulogic;
    signal P0CMDFULL_out : std_ulogic;
    signal P0RDCOUNT_out : std_logic_vector(6 downto 0);
    signal P0RDDATA_out : std_logic_vector(31 downto 0);
    signal P0RDEMPTY_out : std_ulogic;
    signal P0RDERROR_out : std_ulogic;
    signal P0RDFULL_out : std_ulogic;
    signal P0RDOVERFLOW_out : std_ulogic;
    signal P0WRCOUNT_out : std_logic_vector(6 downto 0);
    signal P0WREMPTY_out : std_ulogic;
    signal P0WRERROR_out : std_ulogic;
    signal P0WRFULL_out : std_ulogic;
    signal P0WRUNDERRUN_out : std_ulogic;
    signal P1CMDEMPTY_out : std_ulogic;
    signal P1CMDFULL_out : std_ulogic;
    signal P1RDCOUNT_out : std_logic_vector(6 downto 0);
    signal P1RDDATA_out : std_logic_vector(31 downto 0);
    signal P1RDEMPTY_out : std_ulogic;
    signal P1RDERROR_out : std_ulogic;
    signal P1RDFULL_out : std_ulogic;
    signal P1RDOVERFLOW_out : std_ulogic;
    signal P1WRCOUNT_out : std_logic_vector(6 downto 0);
    signal P1WREMPTY_out : std_ulogic;
    signal P1WRERROR_out : std_ulogic;
    signal P1WRFULL_out : std_ulogic;
    signal P1WRUNDERRUN_out : std_ulogic;
    signal P2CMDEMPTY_out : std_ulogic;
    signal P2CMDFULL_out : std_ulogic;
    signal P2COUNT_out : std_logic_vector(6 downto 0);
    signal P2EMPTY_out : std_ulogic;
    signal P2ERROR_out : std_ulogic;
    signal P2FULL_out : std_ulogic;
    signal P2RDDATA_out : std_logic_vector(31 downto 0);
    signal P2RDOVERFLOW_out : std_ulogic;
    signal P2WRUNDERRUN_out : std_ulogic;
    signal P3CMDEMPTY_out : std_ulogic;
    signal P3CMDFULL_out : std_ulogic;
    signal P3COUNT_out : std_logic_vector(6 downto 0);
    signal P3EMPTY_out : std_ulogic;
    signal P3ERROR_out : std_ulogic;
    signal P3FULL_out : std_ulogic;
    signal P3RDDATA_out : std_logic_vector(31 downto 0);
    signal P3RDOVERFLOW_out : std_ulogic;
    signal P3WRUNDERRUN_out : std_ulogic;
    signal P4CMDEMPTY_out : std_ulogic;
    signal P4CMDFULL_out : std_ulogic;
    signal P4COUNT_out : std_logic_vector(6 downto 0);
    signal P4EMPTY_out : std_ulogic;
    signal P4ERROR_out : std_ulogic;
    signal P4FULL_out : std_ulogic;
    signal P4RDDATA_out : std_logic_vector(31 downto 0);
    signal P4RDOVERFLOW_out : std_ulogic;
    signal P4WRUNDERRUN_out : std_ulogic;
    signal P5CMDEMPTY_out : std_ulogic;
    signal P5CMDFULL_out : std_ulogic;
    signal P5COUNT_out : std_logic_vector(6 downto 0);
    signal P5EMPTY_out : std_ulogic;
    signal P5ERROR_out : std_ulogic;
    signal P5FULL_out : std_ulogic;
    signal P5RDDATA_out : std_logic_vector(31 downto 0);
    signal P5RDOVERFLOW_out : std_ulogic;
    signal P5WRUNDERRUN_out : std_ulogic;
    signal RAS_out : std_ulogic;
    signal RST_out : std_ulogic;
    signal SELFREFRESHMODE_out : std_ulogic;
    signal STATUS_out : std_logic_vector(31 downto 0);
    signal UDMN_out : std_ulogic;
    signal UDMP_out : std_ulogic;
    signal UOCALSTART_out : std_ulogic;
    signal UOCMDREADYIN_out : std_ulogic;
    signal UODATAVALID_out : std_ulogic;
    signal UODATA_out : std_logic_vector(7 downto 0);
    signal UODONECAL_out : std_ulogic;
    signal UOREFRSHFLAG_out : std_ulogic;
    signal UOSDO_out : std_ulogic;
    signal WE_out : std_ulogic;
    
    signal ADDR_outdelay : std_logic_vector(14 downto 0);
    signal BA_outdelay : std_logic_vector(2 downto 0);
    signal CAS_outdelay : std_ulogic;
    signal CKE_outdelay : std_ulogic;
    signal DQIOWEN0_outdelay : std_ulogic;
    signal DQON_outdelay : std_logic_vector(15 downto 0);
    signal DQOP_outdelay : std_logic_vector(15 downto 0);
    signal DQSIOWEN90N_outdelay : std_ulogic;
    signal DQSIOWEN90P_outdelay : std_ulogic;
    signal IOIDRPADDR_outdelay : std_logic_vector(4 downto 0);
    signal IOIDRPADD_outdelay : std_ulogic;
    signal IOIDRPBROADCAST_outdelay : std_ulogic;
    signal IOIDRPCLK_outdelay : std_ulogic;
    signal IOIDRPCS_outdelay : std_ulogic;
    signal IOIDRPSDO_outdelay : std_ulogic;
    signal IOIDRPTRAIN_outdelay : std_ulogic;
    signal IOIDRPUPDATE_outdelay : std_ulogic;
    signal LDMN_outdelay : std_ulogic;
    signal LDMP_outdelay : std_ulogic;
    signal ODT_outdelay : std_ulogic;
    signal P0CMDEMPTY_outdelay : std_ulogic;
    signal P0CMDFULL_outdelay : std_ulogic;
    signal P0RDCOUNT_outdelay : std_logic_vector(6 downto 0);
    signal P0RDDATA_outdelay : std_logic_vector(31 downto 0);
    signal P0RDEMPTY_outdelay : std_ulogic;
    signal P0RDERROR_outdelay : std_ulogic;
    signal P0RDFULL_outdelay : std_ulogic;
    signal P0RDOVERFLOW_outdelay : std_ulogic;
    signal P0WRCOUNT_outdelay : std_logic_vector(6 downto 0);
    signal P0WREMPTY_outdelay : std_ulogic;
    signal P0WRERROR_outdelay : std_ulogic;
    signal P0WRFULL_outdelay : std_ulogic;
    signal P0WRUNDERRUN_outdelay : std_ulogic;
    signal P1CMDEMPTY_outdelay : std_ulogic;
    signal P1CMDFULL_outdelay : std_ulogic;
    signal P1RDCOUNT_outdelay : std_logic_vector(6 downto 0);
    signal P1RDDATA_outdelay : std_logic_vector(31 downto 0);
    signal P1RDEMPTY_outdelay : std_ulogic;
    signal P1RDERROR_outdelay : std_ulogic;
    signal P1RDFULL_outdelay : std_ulogic;
    signal P1RDOVERFLOW_outdelay : std_ulogic;
    signal P1WRCOUNT_outdelay : std_logic_vector(6 downto 0);
    signal P1WREMPTY_outdelay : std_ulogic;
    signal P1WRERROR_outdelay : std_ulogic;
    signal P1WRFULL_outdelay : std_ulogic;
    signal P1WRUNDERRUN_outdelay : std_ulogic;
    signal P2CMDEMPTY_outdelay : std_ulogic;
    signal P2CMDFULL_outdelay : std_ulogic;
    signal P2COUNT_outdelay : std_logic_vector(6 downto 0);
    signal P2EMPTY_outdelay : std_ulogic;
    signal P2ERROR_outdelay : std_ulogic;
    signal P2FULL_outdelay : std_ulogic;
    signal P2RDDATA_outdelay : std_logic_vector(31 downto 0);
    signal P2RDOVERFLOW_outdelay : std_ulogic;
    signal P2WRUNDERRUN_outdelay : std_ulogic;
    signal P3CMDEMPTY_outdelay : std_ulogic;
    signal P3CMDFULL_outdelay : std_ulogic;
    signal P3COUNT_outdelay : std_logic_vector(6 downto 0);
    signal P3EMPTY_outdelay : std_ulogic;
    signal P3ERROR_outdelay : std_ulogic;
    signal P3FULL_outdelay : std_ulogic;
    signal P3RDDATA_outdelay : std_logic_vector(31 downto 0);
    signal P3RDOVERFLOW_outdelay : std_ulogic;
    signal P3WRUNDERRUN_outdelay : std_ulogic;
    signal P4CMDEMPTY_outdelay : std_ulogic;
    signal P4CMDFULL_outdelay : std_ulogic;
    signal P4COUNT_outdelay : std_logic_vector(6 downto 0);
    signal P4EMPTY_outdelay : std_ulogic;
    signal P4ERROR_outdelay : std_ulogic;
    signal P4FULL_outdelay : std_ulogic;
    signal P4RDDATA_outdelay : std_logic_vector(31 downto 0);
    signal P4RDOVERFLOW_outdelay : std_ulogic;
    signal P4WRUNDERRUN_outdelay : std_ulogic;
    signal P5CMDEMPTY_outdelay : std_ulogic;
    signal P5CMDFULL_outdelay : std_ulogic;
    signal P5COUNT_outdelay : std_logic_vector(6 downto 0);
    signal P5EMPTY_outdelay : std_ulogic;
    signal P5ERROR_outdelay : std_ulogic;
    signal P5FULL_outdelay : std_ulogic;
    signal P5RDDATA_outdelay : std_logic_vector(31 downto 0);
    signal P5RDOVERFLOW_outdelay : std_ulogic;
    signal P5WRUNDERRUN_outdelay : std_ulogic;
    signal RAS_outdelay : std_ulogic;
    signal RST_outdelay : std_ulogic;
    signal SELFREFRESHMODE_outdelay : std_ulogic;
    signal STATUS_outdelay : std_logic_vector(31 downto 0);
    signal UDMN_outdelay : std_ulogic;
    signal UDMP_outdelay : std_ulogic;
    signal UOCALSTART_outdelay : std_ulogic;
    signal UOCMDREADYIN_outdelay : std_ulogic;
    signal UODATAVALID_outdelay : std_ulogic;
    signal UODATA_outdelay : std_logic_vector(7 downto 0);
    signal UODONECAL_outdelay : std_ulogic;
    signal UOREFRSHFLAG_outdelay : std_ulogic;
    signal UOSDO_outdelay : std_ulogic;
    signal WE_outdelay : std_ulogic;
    
    signal DQI_ipd : std_logic_vector(15 downto 0);
    signal DQSIOIN_ipd : std_ulogic;
    signal DQSIOIP_ipd : std_ulogic;
    signal IOIDRPSDI_ipd : std_ulogic;
    signal P0ARBEN_ipd : std_ulogic;
    signal P0CMDBA_ipd : std_logic_vector(2 downto 0);
    signal P0CMDBL_ipd : std_logic_vector(5 downto 0);
    signal P0CMDCA_ipd : std_logic_vector(11 downto 0);
    signal P0CMDCLK_ipd : std_ulogic;
    signal P0CMDEN_ipd : std_ulogic;
    signal P0CMDINSTR_ipd : std_logic_vector(2 downto 0);
    signal P0CMDRA_ipd : std_logic_vector(14 downto 0);
    signal P0RDCLK_ipd : std_ulogic;
    signal P0RDEN_ipd : std_ulogic;
    signal P0RWRMASK_ipd : std_logic_vector(3 downto 0);
    signal P0WRCLK_ipd : std_ulogic;
    signal P0WRDATA_ipd : std_logic_vector(31 downto 0);
    signal P0WREN_ipd : std_ulogic;
    signal P1ARBEN_ipd : std_ulogic;
    signal P1CMDBA_ipd : std_logic_vector(2 downto 0);
    signal P1CMDBL_ipd : std_logic_vector(5 downto 0);
    signal P1CMDCA_ipd : std_logic_vector(11 downto 0);
    signal P1CMDCLK_ipd : std_ulogic;
    signal P1CMDEN_ipd : std_ulogic;
    signal P1CMDINSTR_ipd : std_logic_vector(2 downto 0);
    signal P1CMDRA_ipd : std_logic_vector(14 downto 0);
    signal P1RDCLK_ipd : std_ulogic;
    signal P1RDEN_ipd : std_ulogic;
    signal P1RWRMASK_ipd : std_logic_vector(3 downto 0);
    signal P1WRCLK_ipd : std_ulogic;
    signal P1WRDATA_ipd : std_logic_vector(31 downto 0);
    signal P1WREN_ipd : std_ulogic;
    signal P2ARBEN_ipd : std_ulogic;
    signal P2CLK_ipd : std_ulogic;
    signal P2CMDBA_ipd : std_logic_vector(2 downto 0);
    signal P2CMDBL_ipd : std_logic_vector(5 downto 0);
    signal P2CMDCA_ipd : std_logic_vector(11 downto 0);
    signal P2CMDCLK_ipd : std_ulogic;
    signal P2CMDEN_ipd : std_ulogic;
    signal P2CMDINSTR_ipd : std_logic_vector(2 downto 0);
    signal P2CMDRA_ipd : std_logic_vector(14 downto 0);
    signal P2EN_ipd : std_ulogic;
    signal P2WRDATA_ipd : std_logic_vector(31 downto 0);
    signal P2WRMASK_ipd : std_logic_vector(3 downto 0);
    signal P3ARBEN_ipd : std_ulogic;
    signal P3CLK_ipd : std_ulogic;
    signal P3CMDBA_ipd : std_logic_vector(2 downto 0);
    signal P3CMDBL_ipd : std_logic_vector(5 downto 0);
    signal P3CMDCA_ipd : std_logic_vector(11 downto 0);
    signal P3CMDCLK_ipd : std_ulogic;
    signal P3CMDEN_ipd : std_ulogic;
    signal P3CMDINSTR_ipd : std_logic_vector(2 downto 0);
    signal P3CMDRA_ipd : std_logic_vector(14 downto 0);
    signal P3EN_ipd : std_ulogic;
    signal P3WRDATA_ipd : std_logic_vector(31 downto 0);
    signal P3WRMASK_ipd : std_logic_vector(3 downto 0);
    signal P4ARBEN_ipd : std_ulogic;
    signal P4CLK_ipd : std_ulogic;
    signal P4CMDBA_ipd : std_logic_vector(2 downto 0);
    signal P4CMDBL_ipd : std_logic_vector(5 downto 0);
    signal P4CMDCA_ipd : std_logic_vector(11 downto 0);
    signal P4CMDCLK_ipd : std_ulogic;
    signal P4CMDEN_ipd : std_ulogic;
    signal P4CMDINSTR_ipd : std_logic_vector(2 downto 0);
    signal P4CMDRA_ipd : std_logic_vector(14 downto 0);
    signal P4EN_ipd : std_ulogic;
    signal P4WRDATA_ipd : std_logic_vector(31 downto 0);
    signal P4WRMASK_ipd : std_logic_vector(3 downto 0);
    signal P5ARBEN_ipd : std_ulogic;
    signal P5CLK_ipd : std_ulogic;
    signal P5CMDBA_ipd : std_logic_vector(2 downto 0);
    signal P5CMDBL_ipd : std_logic_vector(5 downto 0);
    signal P5CMDCA_ipd : std_logic_vector(11 downto 0);
    signal P5CMDCLK_ipd : std_ulogic;
    signal P5CMDEN_ipd : std_ulogic;
    signal P5CMDINSTR_ipd : std_logic_vector(2 downto 0);
    signal P5CMDRA_ipd : std_logic_vector(14 downto 0);
    signal P5EN_ipd : std_ulogic;
    signal P5WRDATA_ipd : std_logic_vector(31 downto 0);
    signal P5WRMASK_ipd : std_logic_vector(3 downto 0);
    signal PLLCE_ipd : std_logic_vector(1 downto 0);
    signal PLLCLK_ipd : std_logic_vector(1 downto 0);
    signal PLLLOCK_ipd : std_ulogic;
    signal RECAL_ipd : std_ulogic;
    signal SELFREFRESHENTER_ipd : std_ulogic;
    signal SYSRST_ipd : std_ulogic;
    signal UDQSIOIN_ipd : std_ulogic;
    signal UDQSIOIP_ipd : std_ulogic;
    signal UIADDR_ipd : std_logic_vector(4 downto 0);
    signal UIADD_ipd : std_ulogic;
    signal UIBROADCAST_ipd : std_ulogic;
    signal UICLK_ipd : std_ulogic;
    signal UICMDEN_ipd : std_ulogic;
    signal UICMDIN_ipd : std_ulogic;
    signal UICMD_ipd : std_ulogic;
    signal UICS_ipd : std_ulogic;
    signal UIDONECAL_ipd : std_ulogic;
    signal UIDQCOUNT_ipd : std_logic_vector(3 downto 0);
    signal UIDQLOWERDEC_ipd : std_ulogic;
    signal UIDQLOWERINC_ipd : std_ulogic;
    signal UIDQUPPERDEC_ipd : std_ulogic;
    signal UIDQUPPERINC_ipd : std_ulogic;
    signal UIDRPUPDATE_ipd : std_ulogic;
    signal UILDQSDEC_ipd : std_ulogic;
    signal UILDQSINC_ipd : std_ulogic;
    signal UIREAD_ipd : std_ulogic;
    signal UISDI_ipd : std_ulogic;
    signal UIUDQSDEC_ipd : std_ulogic;
    signal UIUDQSINC_ipd : std_ulogic;
    
    signal IOIDRPSDI_UICLK_dly : std_ulogic;
    signal P0ARBEN_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal P0CMDBA_P0CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P0CMDBL_P0CMDCLK_dly : std_logic_vector(5 downto 0);
    signal P0CMDCA_P0CMDCLK_dly : std_logic_vector(11 downto 0);
    signal P0CMDCLK_dly : std_ulogic;
    signal P0CMDEN_P0CMDCLK_dly : std_ulogic;
    signal P0CMDINSTR_P0CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P0CMDRA_P0CMDCLK_dly : std_logic_vector(14 downto 0);
    signal P0RDCLK_dly : std_ulogic;
    signal P0RDEN_P0RDCLK_dly : std_ulogic;
    signal P0RWRMASK_P0WRCLK_dly : std_logic_vector(3 downto 0);
    signal P0WRCLK_dly : std_ulogic;
    signal P0WRDATA_P0WRCLK_dly : std_logic_vector(31 downto 0);
    signal P0WREN_P0WRCLK_dly : std_ulogic;
    signal P1ARBEN_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal P1CMDBA_P1CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P1CMDBL_P1CMDCLK_dly : std_logic_vector(5 downto 0);
    signal P1CMDCA_P1CMDCLK_dly : std_logic_vector(11 downto 0);
    signal P1CMDCLK_dly : std_ulogic;
    signal P1CMDEN_P1CMDCLK_dly : std_ulogic;
    signal P1CMDINSTR_P1CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P1CMDRA_P1CMDCLK_dly : std_logic_vector(14 downto 0);
    signal P1RDCLK_dly : std_ulogic;
    signal P1RDEN_P1RDCLK_dly : std_ulogic;
    signal P1RWRMASK_P1WRCLK_dly : std_logic_vector(3 downto 0);
    signal P1WRCLK_dly : std_ulogic;
    signal P1WRDATA_P1WRCLK_dly : std_logic_vector(31 downto 0);
    signal P1WREN_P1WRCLK_dly : std_ulogic;
    signal P2ARBEN_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal P2CLK_dly : std_ulogic;
    signal P2CMDBA_P2CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P2CMDBL_P2CMDCLK_dly : std_logic_vector(5 downto 0);
    signal P2CMDCA_P2CMDCLK_dly : std_logic_vector(11 downto 0);
    signal P2CMDCLK_dly : std_ulogic;
    signal P2CMDEN_P2CMDCLK_dly : std_ulogic;
    signal P2CMDINSTR_P2CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P2CMDRA_P2CMDCLK_dly : std_logic_vector(14 downto 0);
    signal P2EN_P2CLK_dly : std_ulogic;
    signal P2WRDATA_P2CLK_dly : std_logic_vector(31 downto 0);
    signal P2WRMASK_P2CLK_dly : std_logic_vector(3 downto 0);
    signal P3ARBEN_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal P3CLK_dly : std_ulogic;
    signal P3CMDBA_P3CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P3CMDBL_P3CMDCLK_dly : std_logic_vector(5 downto 0);
    signal P3CMDCA_P3CMDCLK_dly : std_logic_vector(11 downto 0);
    signal P3CMDCLK_dly : std_ulogic;
    signal P3CMDEN_P3CMDCLK_dly : std_ulogic;
    signal P3CMDINSTR_P3CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P3CMDRA_P3CMDCLK_dly : std_logic_vector(14 downto 0);
    signal P3EN_P3CLK_dly : std_ulogic;
    signal P3WRDATA_P3CLK_dly : std_logic_vector(31 downto 0);
    signal P3WRMASK_P3CLK_dly : std_logic_vector(3 downto 0);
    signal P4ARBEN_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal P4CLK_dly : std_ulogic;
    signal P4CMDBA_P4CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P4CMDBL_P4CMDCLK_dly : std_logic_vector(5 downto 0);
    signal P4CMDCA_P4CMDCLK_dly : std_logic_vector(11 downto 0);
    signal P4CMDCLK_dly : std_ulogic;
    signal P4CMDEN_P4CMDCLK_dly : std_ulogic;
    signal P4CMDINSTR_P4CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P4CMDRA_P4CMDCLK_dly : std_logic_vector(14 downto 0);
    signal P4EN_P4CLK_dly : std_ulogic;
    signal P4WRDATA_P4CLK_dly : std_logic_vector(31 downto 0);
    signal P4WRMASK_P4CLK_dly : std_logic_vector(3 downto 0);
    signal P5ARBEN_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal P5CLK_dly : std_ulogic;
    signal P5CMDBA_P5CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P5CMDBL_P5CMDCLK_dly : std_logic_vector(5 downto 0);
    signal P5CMDCA_P5CMDCLK_dly : std_logic_vector(11 downto 0);
    signal P5CMDCLK_dly : std_ulogic;
    signal P5CMDEN_P5CMDCLK_dly : std_ulogic;
    signal P5CMDINSTR_P5CMDCLK_dly : std_logic_vector(2 downto 0);
    signal P5CMDRA_P5CMDCLK_dly : std_logic_vector(14 downto 0);
    signal P5EN_P5CLK_dly : std_ulogic;
    signal P5WRDATA_P5CLK_dly : std_logic_vector(31 downto 0);
    signal P5WRMASK_P5CLK_dly : std_logic_vector(3 downto 0);
    signal PLLCE_PLLCLK_dly : std_logic_vector(3 downto 0);
    signal PLLCLK_dly : std_logic_vector(1 downto 0);
    signal PLLLOCK_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal RECAL_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal SELFREFRESHENTER_PLLCLK_dly : std_logic_vector(1 downto 0);
    signal SYSRST_dly : std_ulogic;
    signal UIADDR_UICLK_dly : std_logic_vector(4 downto 0);
    signal UIADD_UICLK_dly : std_ulogic;
    signal UIBROADCAST_UICLK_dly : std_ulogic;
    signal UICLK_dly : std_ulogic;
    signal UICMDEN_UICLK_dly : std_ulogic;
    signal UICMDIN_UICLK_dly : std_ulogic;
    signal UICMD_UICLK_dly : std_ulogic;
    signal UICS_UICLK_dly : std_ulogic;
    signal UIDONECAL_UICLK_dly : std_ulogic;
    signal UIDQCOUNT_UICLK_dly : std_logic_vector(3 downto 0);
    signal UIDQLOWERDEC_UICLK_dly : std_ulogic;
    signal UIDQLOWERINC_UICLK_dly : std_ulogic;
    signal UIDQUPPERDEC_UICLK_dly : std_ulogic;
    signal UIDQUPPERINC_UICLK_dly : std_ulogic;
    signal UIDRPUPDATE_UICLK_dly : std_ulogic;
    signal UILDQSDEC_UICLK_dly : std_ulogic;
    signal UILDQSINC_UICLK_dly : std_ulogic;
    signal UIREAD_UICLK_dly : std_ulogic;
    signal UISDI_UICLK_dly : std_ulogic;
    signal UIUDQSDEC_UICLK_dly : std_ulogic;
    signal UIUDQSINC_UICLK_dly : std_ulogic;
    
    signal DQI_indelay : std_logic_vector(15 downto 0);
    signal DQSIOIN_indelay : std_ulogic;
    signal DQSIOIP_indelay : std_ulogic;
    signal IOIDRPSDI_indelay : std_ulogic;
    signal P0ARBEN_indelay : std_ulogic;
    signal P0CMDBA_indelay : std_logic_vector(2 downto 0);
    signal P0CMDBL_indelay : std_logic_vector(5 downto 0);
    signal P0CMDCA_indelay : std_logic_vector(11 downto 0);
    signal P0CMDCLK_indelay : std_ulogic;
    signal P0CMDEN_indelay : std_ulogic;
    signal P0CMDINSTR_indelay : std_logic_vector(2 downto 0);
    signal P0CMDRA_indelay : std_logic_vector(14 downto 0);
    signal P0RDCLK_indelay : std_ulogic;
    signal P0RDEN_indelay : std_ulogic;
    signal P0RWRMASK_indelay : std_logic_vector(3 downto 0);
    signal P0WRCLK_indelay : std_ulogic;
    signal P0WRDATA_indelay : std_logic_vector(31 downto 0);
    signal P0WREN_indelay : std_ulogic;
    signal P1ARBEN_indelay : std_ulogic;
    signal P1CMDBA_indelay : std_logic_vector(2 downto 0);
    signal P1CMDBL_indelay : std_logic_vector(5 downto 0);
    signal P1CMDCA_indelay : std_logic_vector(11 downto 0);
    signal P1CMDCLK_indelay : std_ulogic;
    signal P1CMDEN_indelay : std_ulogic;
    signal P1CMDINSTR_indelay : std_logic_vector(2 downto 0);
    signal P1CMDRA_indelay : std_logic_vector(14 downto 0);
    signal P1RDCLK_indelay : std_ulogic;
    signal P1RDEN_indelay : std_ulogic;
    signal P1RWRMASK_indelay : std_logic_vector(3 downto 0);
    signal P1WRCLK_indelay : std_ulogic;
    signal P1WRDATA_indelay : std_logic_vector(31 downto 0);
    signal P1WREN_indelay : std_ulogic;
    signal P2ARBEN_indelay : std_ulogic;
    signal P2CLK_indelay : std_ulogic;
    signal P2CMDBA_indelay : std_logic_vector(2 downto 0);
    signal P2CMDBL_indelay : std_logic_vector(5 downto 0);
    signal P2CMDCA_indelay : std_logic_vector(11 downto 0);
    signal P2CMDCLK_indelay : std_ulogic;
    signal P2CMDEN_indelay : std_ulogic;
    signal P2CMDINSTR_indelay : std_logic_vector(2 downto 0);
    signal P2CMDRA_indelay : std_logic_vector(14 downto 0);
    signal P2EN_indelay : std_ulogic;
    signal P2WRDATA_indelay : std_logic_vector(31 downto 0);
    signal P2WRMASK_indelay : std_logic_vector(3 downto 0);
    signal P3ARBEN_indelay : std_ulogic;
    signal P3CLK_indelay : std_ulogic;
    signal P3CMDBA_indelay : std_logic_vector(2 downto 0);
    signal P3CMDBL_indelay : std_logic_vector(5 downto 0);
    signal P3CMDCA_indelay : std_logic_vector(11 downto 0);
    signal P3CMDCLK_indelay : std_ulogic;
    signal P3CMDEN_indelay : std_ulogic;
    signal P3CMDINSTR_indelay : std_logic_vector(2 downto 0);
    signal P3CMDRA_indelay : std_logic_vector(14 downto 0);
    signal P3EN_indelay : std_ulogic;
    signal P3WRDATA_indelay : std_logic_vector(31 downto 0);
    signal P3WRMASK_indelay : std_logic_vector(3 downto 0);
    signal P4ARBEN_indelay : std_ulogic;
    signal P4CLK_indelay : std_ulogic;
    signal P4CMDBA_indelay : std_logic_vector(2 downto 0);
    signal P4CMDBL_indelay : std_logic_vector(5 downto 0);
    signal P4CMDCA_indelay : std_logic_vector(11 downto 0);
    signal P4CMDCLK_indelay : std_ulogic;
    signal P4CMDEN_indelay : std_ulogic;
    signal P4CMDINSTR_indelay : std_logic_vector(2 downto 0);
    signal P4CMDRA_indelay : std_logic_vector(14 downto 0);
    signal P4EN_indelay : std_ulogic;
    signal P4WRDATA_indelay : std_logic_vector(31 downto 0);
    signal P4WRMASK_indelay : std_logic_vector(3 downto 0);
    signal P5ARBEN_indelay : std_ulogic;
    signal P5CLK_indelay : std_ulogic;
    signal P5CMDBA_indelay : std_logic_vector(2 downto 0);
    signal P5CMDBL_indelay : std_logic_vector(5 downto 0);
    signal P5CMDCA_indelay : std_logic_vector(11 downto 0);
    signal P5CMDCLK_indelay : std_ulogic;
    signal P5CMDEN_indelay : std_ulogic;
    signal P5CMDINSTR_indelay : std_logic_vector(2 downto 0);
    signal P5CMDRA_indelay : std_logic_vector(14 downto 0);
    signal P5EN_indelay : std_ulogic;
    signal P5WRDATA_indelay : std_logic_vector(31 downto 0);
    signal P5WRMASK_indelay : std_logic_vector(3 downto 0);
    signal PLLCE_indelay : std_logic_vector(1 downto 0);
    signal PLLCLK_indelay : std_logic_vector(1 downto 0);
    signal PLLLOCK_indelay : std_ulogic;
    signal RECAL_indelay : std_ulogic;
    signal SELFREFRESHENTER_indelay : std_ulogic;
    signal SYSRST_indelay : std_ulogic;
    signal UDQSIOIN_indelay : std_ulogic;
    signal UDQSIOIP_indelay : std_ulogic;
    signal UIADDR_indelay : std_logic_vector(4 downto 0);
    signal UIADD_indelay : std_ulogic;
    signal UIBROADCAST_indelay : std_ulogic;
    signal UICLK_indelay : std_ulogic;
    signal UICMDEN_indelay : std_ulogic;
    signal UICMDIN_indelay : std_ulogic;
    signal UICMD_indelay : std_ulogic;
    signal UICS_indelay : std_ulogic;
    signal UIDONECAL_indelay : std_ulogic;
    signal UIDQCOUNT_indelay : std_logic_vector(3 downto 0);
    signal UIDQLOWERDEC_indelay : std_ulogic;
    signal UIDQLOWERINC_indelay : std_ulogic;
    signal UIDQUPPERDEC_indelay : std_ulogic;
    signal UIDQUPPERINC_indelay : std_ulogic;
    signal UIDRPUPDATE_indelay : std_ulogic;
    signal UILDQSDEC_indelay : std_ulogic;
    signal UILDQSINC_indelay : std_ulogic;
    signal UIREAD_indelay : std_ulogic;
    signal UISDI_indelay : std_ulogic;
    signal UIUDQSDEC_indelay : std_ulogic;
    signal UIUDQSINC_indelay : std_ulogic;
    
    signal DQI_indly : std_logic_vector(15 downto 0);
    signal DQSIOIN_indly : std_ulogic;
    signal DQSIOIP_indly : std_ulogic;
    signal IOIDRPSDI_indly : std_ulogic;
    signal P0ARBEN_indly : std_ulogic;
    signal P0CMDBA_indly : std_logic_vector(2 downto 0);
    signal P0CMDBL_indly : std_logic_vector(5 downto 0);
    signal P0CMDCA_indly : std_logic_vector(11 downto 0);
    signal P0CMDCLK_indly : std_ulogic;
    signal P0CMDEN_indly : std_ulogic;
    signal P0CMDINSTR_indly : std_logic_vector(2 downto 0);
    signal P0CMDRA_indly : std_logic_vector(14 downto 0);
    signal P0RDCLK_indly : std_ulogic;
    signal P0RDEN_indly : std_ulogic;
    signal P0RWRMASK_indly : std_logic_vector(3 downto 0);
    signal P0WRCLK_indly : std_ulogic;
    signal P0WRDATA_indly : std_logic_vector(31 downto 0);
    signal P0WREN_indly : std_ulogic;
    signal P1ARBEN_indly : std_ulogic;
    signal P1CMDBA_indly : std_logic_vector(2 downto 0);
    signal P1CMDBL_indly : std_logic_vector(5 downto 0);
    signal P1CMDCA_indly : std_logic_vector(11 downto 0);
    signal P1CMDCLK_indly : std_ulogic;
    signal P1CMDEN_indly : std_ulogic;
    signal P1CMDINSTR_indly : std_logic_vector(2 downto 0);
    signal P1CMDRA_indly : std_logic_vector(14 downto 0);
    signal P1RDCLK_indly : std_ulogic;
    signal P1RDEN_indly : std_ulogic;
    signal P1RWRMASK_indly : std_logic_vector(3 downto 0);
    signal P1WRCLK_indly : std_ulogic;
    signal P1WRDATA_indly : std_logic_vector(31 downto 0);
    signal P1WREN_indly : std_ulogic;
    signal P2ARBEN_indly : std_ulogic;
    signal P2CLK_indly : std_ulogic;
    signal P2CMDBA_indly : std_logic_vector(2 downto 0);
    signal P2CMDBL_indly : std_logic_vector(5 downto 0);
    signal P2CMDCA_indly : std_logic_vector(11 downto 0);
    signal P2CMDCLK_indly : std_ulogic;
    signal P2CMDEN_indly : std_ulogic;
    signal P2CMDINSTR_indly : std_logic_vector(2 downto 0);
    signal P2CMDRA_indly : std_logic_vector(14 downto 0);
    signal P2EN_indly : std_ulogic;
    signal P2WRDATA_indly : std_logic_vector(31 downto 0);
    signal P2WRMASK_indly : std_logic_vector(3 downto 0);
    signal P3ARBEN_indly : std_ulogic;
    signal P3CLK_indly : std_ulogic;
    signal P3CMDBA_indly : std_logic_vector(2 downto 0);
    signal P3CMDBL_indly : std_logic_vector(5 downto 0);
    signal P3CMDCA_indly : std_logic_vector(11 downto 0);
    signal P3CMDCLK_indly : std_ulogic;
    signal P3CMDEN_indly : std_ulogic;
    signal P3CMDINSTR_indly : std_logic_vector(2 downto 0);
    signal P3CMDRA_indly : std_logic_vector(14 downto 0);
    signal P3EN_indly : std_ulogic;
    signal P3WRDATA_indly : std_logic_vector(31 downto 0);
    signal P3WRMASK_indly : std_logic_vector(3 downto 0);
    signal P4ARBEN_indly : std_ulogic;
    signal P4CLK_indly : std_ulogic;
    signal P4CMDBA_indly : std_logic_vector(2 downto 0);
    signal P4CMDBL_indly : std_logic_vector(5 downto 0);
    signal P4CMDCA_indly : std_logic_vector(11 downto 0);
    signal P4CMDCLK_indly : std_ulogic;
    signal P4CMDEN_indly : std_ulogic;
    signal P4CMDINSTR_indly : std_logic_vector(2 downto 0);
    signal P4CMDRA_indly : std_logic_vector(14 downto 0);
    signal P4EN_indly : std_ulogic;
    signal P4WRDATA_indly : std_logic_vector(31 downto 0);
    signal P4WRMASK_indly : std_logic_vector(3 downto 0);
    signal P5ARBEN_indly : std_ulogic;
    signal P5CLK_indly : std_ulogic;
    signal P5CMDBA_indly : std_logic_vector(2 downto 0);
    signal P5CMDBL_indly : std_logic_vector(5 downto 0);
    signal P5CMDCA_indly : std_logic_vector(11 downto 0);
    signal P5CMDCLK_indly : std_ulogic;
    signal P5CMDEN_indly : std_ulogic;
    signal P5CMDINSTR_indly : std_logic_vector(2 downto 0);
    signal P5CMDRA_indly : std_logic_vector(14 downto 0);
    signal P5EN_indly : std_ulogic;
    signal P5WRDATA_indly : std_logic_vector(31 downto 0);
    signal P5WRMASK_indly : std_logic_vector(3 downto 0);
    signal PLLCE_indly : std_logic_vector(1 downto 0);
    signal PLLCLK_indly : std_logic_vector(1 downto 0);
    signal PLLLOCK_indly : std_ulogic;
    signal RECAL_indly : std_ulogic;
    signal SELFREFRESHENTER_indly : std_ulogic;
    signal SYSRST_indly : std_ulogic;
    signal UDQSIOIN_indly : std_ulogic;
    signal UDQSIOIP_indly : std_ulogic;
    signal UIADDR_indly : std_logic_vector(4 downto 0);
    signal UIADD_indly : std_ulogic;
    signal UIBROADCAST_indly : std_ulogic;
    signal UICLK_indly : std_ulogic;
    signal UICMDEN_indly : std_ulogic;
    signal UICMDIN_indly : std_ulogic;
    signal UICMD_indly : std_ulogic;
    signal UICS_indly : std_ulogic;
    signal UIDONECAL_indly : std_ulogic;
    signal UIDQCOUNT_indly : std_logic_vector(3 downto 0);
    signal UIDQLOWERDEC_indly : std_ulogic;
    signal UIDQLOWERINC_indly : std_ulogic;
    signal UIDQUPPERDEC_indly : std_ulogic;
    signal UIDQUPPERINC_indly : std_ulogic;
    signal UIDRPUPDATE_indly : std_ulogic;
    signal UILDQSDEC_indly : std_ulogic;
    signal UILDQSINC_indly : std_ulogic;
    signal UIREAD_indly : std_ulogic;
    signal UISDI_indly : std_ulogic;
    signal UIUDQSDEC_indly : std_ulogic;
    signal UIUDQSINC_indly : std_ulogic;

-- <!--Aldec correction start
	signal GSR_local : std_ulogic;
-- Aldec correction end -->
    
   signal PLLCLK_0 : std_ulogic ;
   signal PLLCLK_1 : std_ulogic ;
    begin
    
    WireDelay : block
    begin
      DQI_DELAY : for i in 0 to 15 generate
        VitalWireDelay (DQI_ipd(i),DQI(i),tipd_DQI(i));
      end generate DQI_DELAY;
      P0CMDBA_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P0CMDBA_ipd(i),P0CMDBA(i),tipd_P0CMDBA(i));
      end generate P0CMDBA_DELAY;
      P0CMDBL_DELAY : for i in 0 to 5 generate
        VitalWireDelay (P0CMDBL_ipd(i),P0CMDBL(i),tipd_P0CMDBL(i));
      end generate P0CMDBL_DELAY;
      P0CMDCA_DELAY : for i in 0 to 11 generate
        VitalWireDelay (P0CMDCA_ipd(i),P0CMDCA(i),tipd_P0CMDCA(i));
      end generate P0CMDCA_DELAY;
      P0CMDINSTR_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P0CMDINSTR_ipd(i),P0CMDINSTR(i),tipd_P0CMDINSTR(i));
      end generate P0CMDINSTR_DELAY;
      P0CMDRA_DELAY : for i in 0 to 14 generate
        VitalWireDelay (P0CMDRA_ipd(i),P0CMDRA(i),tipd_P0CMDRA(i));
      end generate P0CMDRA_DELAY;
      P0RWRMASK_DELAY : for i in 0 to 3 generate
        VitalWireDelay (P0RWRMASK_ipd(i),P0RWRMASK(i),tipd_P0RWRMASK(i));
      end generate P0RWRMASK_DELAY;
      P0WRDATA_DELAY : for i in 0 to 31 generate
        VitalWireDelay (P0WRDATA_ipd(i),P0WRDATA(i),tipd_P0WRDATA(i));
      end generate P0WRDATA_DELAY;
      P1CMDBA_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P1CMDBA_ipd(i),P1CMDBA(i),tipd_P1CMDBA(i));
      end generate P1CMDBA_DELAY;
      P1CMDBL_DELAY : for i in 0 to 5 generate
        VitalWireDelay (P1CMDBL_ipd(i),P1CMDBL(i),tipd_P1CMDBL(i));
      end generate P1CMDBL_DELAY;
      P1CMDCA_DELAY : for i in 0 to 11 generate
        VitalWireDelay (P1CMDCA_ipd(i),P1CMDCA(i),tipd_P1CMDCA(i));
      end generate P1CMDCA_DELAY;
      P1CMDINSTR_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P1CMDINSTR_ipd(i),P1CMDINSTR(i),tipd_P1CMDINSTR(i));
      end generate P1CMDINSTR_DELAY;
      P1CMDRA_DELAY : for i in 0 to 14 generate
        VitalWireDelay (P1CMDRA_ipd(i),P1CMDRA(i),tipd_P1CMDRA(i));
      end generate P1CMDRA_DELAY;
      P1RWRMASK_DELAY : for i in 0 to 3 generate
        VitalWireDelay (P1RWRMASK_ipd(i),P1RWRMASK(i),tipd_P1RWRMASK(i));
      end generate P1RWRMASK_DELAY;
      P1WRDATA_DELAY : for i in 0 to 31 generate
        VitalWireDelay (P1WRDATA_ipd(i),P1WRDATA(i),tipd_P1WRDATA(i));
      end generate P1WRDATA_DELAY;
      P2CMDBA_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P2CMDBA_ipd(i),P2CMDBA(i),tipd_P2CMDBA(i));
      end generate P2CMDBA_DELAY;
      P2CMDBL_DELAY : for i in 0 to 5 generate
        VitalWireDelay (P2CMDBL_ipd(i),P2CMDBL(i),tipd_P2CMDBL(i));
      end generate P2CMDBL_DELAY;
      P2CMDCA_DELAY : for i in 0 to 11 generate
        VitalWireDelay (P2CMDCA_ipd(i),P2CMDCA(i),tipd_P2CMDCA(i));
      end generate P2CMDCA_DELAY;
      P2CMDINSTR_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P2CMDINSTR_ipd(i),P2CMDINSTR(i),tipd_P2CMDINSTR(i));
      end generate P2CMDINSTR_DELAY;
      P2CMDRA_DELAY : for i in 0 to 14 generate
        VitalWireDelay (P2CMDRA_ipd(i),P2CMDRA(i),tipd_P2CMDRA(i));
      end generate P2CMDRA_DELAY;
      P2WRDATA_DELAY : for i in 0 to 31 generate
        VitalWireDelay (P2WRDATA_ipd(i),P2WRDATA(i),tipd_P2WRDATA(i));
      end generate P2WRDATA_DELAY;
      P2WRMASK_DELAY : for i in 0 to 3 generate
        VitalWireDelay (P2WRMASK_ipd(i),P2WRMASK(i),tipd_P2WRMASK(i));
      end generate P2WRMASK_DELAY;
      P3CMDBA_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P3CMDBA_ipd(i),P3CMDBA(i),tipd_P3CMDBA(i));
      end generate P3CMDBA_DELAY;
      P3CMDBL_DELAY : for i in 0 to 5 generate
        VitalWireDelay (P3CMDBL_ipd(i),P3CMDBL(i),tipd_P3CMDBL(i));
      end generate P3CMDBL_DELAY;
      P3CMDCA_DELAY : for i in 0 to 11 generate
        VitalWireDelay (P3CMDCA_ipd(i),P3CMDCA(i),tipd_P3CMDCA(i));
      end generate P3CMDCA_DELAY;
      P3CMDINSTR_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P3CMDINSTR_ipd(i),P3CMDINSTR(i),tipd_P3CMDINSTR(i));
      end generate P3CMDINSTR_DELAY;
      P3CMDRA_DELAY : for i in 0 to 14 generate
        VitalWireDelay (P3CMDRA_ipd(i),P3CMDRA(i),tipd_P3CMDRA(i));
      end generate P3CMDRA_DELAY;
      P3WRDATA_DELAY : for i in 0 to 31 generate
        VitalWireDelay (P3WRDATA_ipd(i),P3WRDATA(i),tipd_P3WRDATA(i));
      end generate P3WRDATA_DELAY;
      P3WRMASK_DELAY : for i in 0 to 3 generate
        VitalWireDelay (P3WRMASK_ipd(i),P3WRMASK(i),tipd_P3WRMASK(i));
      end generate P3WRMASK_DELAY;
      P4CMDBA_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P4CMDBA_ipd(i),P4CMDBA(i),tipd_P4CMDBA(i));
      end generate P4CMDBA_DELAY;
      P4CMDBL_DELAY : for i in 0 to 5 generate
        VitalWireDelay (P4CMDBL_ipd(i),P4CMDBL(i),tipd_P4CMDBL(i));
      end generate P4CMDBL_DELAY;
      P4CMDCA_DELAY : for i in 0 to 11 generate
        VitalWireDelay (P4CMDCA_ipd(i),P4CMDCA(i),tipd_P4CMDCA(i));
      end generate P4CMDCA_DELAY;
      P4CMDINSTR_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P4CMDINSTR_ipd(i),P4CMDINSTR(i),tipd_P4CMDINSTR(i));
      end generate P4CMDINSTR_DELAY;
      P4CMDRA_DELAY : for i in 0 to 14 generate
        VitalWireDelay (P4CMDRA_ipd(i),P4CMDRA(i),tipd_P4CMDRA(i));
      end generate P4CMDRA_DELAY;
      P4WRDATA_DELAY : for i in 0 to 31 generate
        VitalWireDelay (P4WRDATA_ipd(i),P4WRDATA(i),tipd_P4WRDATA(i));
      end generate P4WRDATA_DELAY;
      P4WRMASK_DELAY : for i in 0 to 3 generate
        VitalWireDelay (P4WRMASK_ipd(i),P4WRMASK(i),tipd_P4WRMASK(i));
      end generate P4WRMASK_DELAY;
      P5CMDBA_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P5CMDBA_ipd(i),P5CMDBA(i),tipd_P5CMDBA(i));
      end generate P5CMDBA_DELAY;
      P5CMDBL_DELAY : for i in 0 to 5 generate
        VitalWireDelay (P5CMDBL_ipd(i),P5CMDBL(i),tipd_P5CMDBL(i));
      end generate P5CMDBL_DELAY;
      P5CMDCA_DELAY : for i in 0 to 11 generate
        VitalWireDelay (P5CMDCA_ipd(i),P5CMDCA(i),tipd_P5CMDCA(i));
      end generate P5CMDCA_DELAY;
      P5CMDINSTR_DELAY : for i in 0 to 2 generate
        VitalWireDelay (P5CMDINSTR_ipd(i),P5CMDINSTR(i),tipd_P5CMDINSTR(i));
      end generate P5CMDINSTR_DELAY;
      P5CMDRA_DELAY : for i in 0 to 14 generate
        VitalWireDelay (P5CMDRA_ipd(i),P5CMDRA(i),tipd_P5CMDRA(i));
      end generate P5CMDRA_DELAY;
      P5WRDATA_DELAY : for i in 0 to 31 generate
        VitalWireDelay (P5WRDATA_ipd(i),P5WRDATA(i),tipd_P5WRDATA(i));
      end generate P5WRDATA_DELAY;
      P5WRMASK_DELAY : for i in 0 to 3 generate
        VitalWireDelay (P5WRMASK_ipd(i),P5WRMASK(i),tipd_P5WRMASK(i));
      end generate P5WRMASK_DELAY;
      PLLCE_DELAY : for i in 0 to 1 generate
        VitalWireDelay (PLLCE_ipd(i),PLLCE(i),tipd_PLLCE(i));
      end generate PLLCE_DELAY;
      PLLCLK_DELAY : for i in 0 to 1 generate
        VitalWireDelay (PLLCLK_ipd(i),PLLCLK(i),tipd_PLLCLK(i));
      end generate PLLCLK_DELAY;
      UIADDR_DELAY : for i in 0 to 4 generate
        VitalWireDelay (UIADDR_ipd(i),UIADDR(i),tipd_UIADDR(i));
      end generate UIADDR_DELAY;
      UIDQCOUNT_DELAY : for i in 0 to 3 generate
        VitalWireDelay (UIDQCOUNT_ipd(i),UIDQCOUNT(i),tipd_UIDQCOUNT(i));
      end generate UIDQCOUNT_DELAY;
      VitalWireDelay (DQSIOIN_ipd,DQSIOIN,tipd_DQSIOIN);
      VitalWireDelay (DQSIOIP_ipd,DQSIOIP,tipd_DQSIOIP);
      VitalWireDelay (IOIDRPSDI_ipd,IOIDRPSDI,tipd_IOIDRPSDI);
      VitalWireDelay (P0ARBEN_ipd,P0ARBEN,tipd_P0ARBEN);
      VitalWireDelay (P0CMDCLK_ipd,P0CMDCLK,tipd_P0CMDCLK);
      VitalWireDelay (P0CMDEN_ipd,P0CMDEN,tipd_P0CMDEN);
      VitalWireDelay (P0RDCLK_ipd,P0RDCLK,tipd_P0RDCLK);
      VitalWireDelay (P0RDEN_ipd,P0RDEN,tipd_P0RDEN);
      VitalWireDelay (P0WRCLK_ipd,P0WRCLK,tipd_P0WRCLK);
      VitalWireDelay (P0WREN_ipd,P0WREN,tipd_P0WREN);
      VitalWireDelay (P1ARBEN_ipd,P1ARBEN,tipd_P1ARBEN);
      VitalWireDelay (P1CMDCLK_ipd,P1CMDCLK,tipd_P1CMDCLK);
      VitalWireDelay (P1CMDEN_ipd,P1CMDEN,tipd_P1CMDEN);
      VitalWireDelay (P1RDCLK_ipd,P1RDCLK,tipd_P1RDCLK);
      VitalWireDelay (P1RDEN_ipd,P1RDEN,tipd_P1RDEN);
      VitalWireDelay (P1WRCLK_ipd,P1WRCLK,tipd_P1WRCLK);
      VitalWireDelay (P1WREN_ipd,P1WREN,tipd_P1WREN);
      VitalWireDelay (P2ARBEN_ipd,P2ARBEN,tipd_P2ARBEN);
      VitalWireDelay (P2CLK_ipd,P2CLK,tipd_P2CLK);
      VitalWireDelay (P2CMDCLK_ipd,P2CMDCLK,tipd_P2CMDCLK);
      VitalWireDelay (P2CMDEN_ipd,P2CMDEN,tipd_P2CMDEN);
      VitalWireDelay (P2EN_ipd,P2EN,tipd_P2EN);
      VitalWireDelay (P3ARBEN_ipd,P3ARBEN,tipd_P3ARBEN);
      VitalWireDelay (P3CLK_ipd,P3CLK,tipd_P3CLK);
      VitalWireDelay (P3CMDCLK_ipd,P3CMDCLK,tipd_P3CMDCLK);
      VitalWireDelay (P3CMDEN_ipd,P3CMDEN,tipd_P3CMDEN);
      VitalWireDelay (P3EN_ipd,P3EN,tipd_P3EN);
      VitalWireDelay (P4ARBEN_ipd,P4ARBEN,tipd_P4ARBEN);
      VitalWireDelay (P4CLK_ipd,P4CLK,tipd_P4CLK);
      VitalWireDelay (P4CMDCLK_ipd,P4CMDCLK,tipd_P4CMDCLK);
      VitalWireDelay (P4CMDEN_ipd,P4CMDEN,tipd_P4CMDEN);
      VitalWireDelay (P4EN_ipd,P4EN,tipd_P4EN);
      VitalWireDelay (P5ARBEN_ipd,P5ARBEN,tipd_P5ARBEN);
      VitalWireDelay (P5CLK_ipd,P5CLK,tipd_P5CLK);
      VitalWireDelay (P5CMDCLK_ipd,P5CMDCLK,tipd_P5CMDCLK);
      VitalWireDelay (P5CMDEN_ipd,P5CMDEN,tipd_P5CMDEN);
      VitalWireDelay (P5EN_ipd,P5EN,tipd_P5EN);
      VitalWireDelay (PLLLOCK_ipd,PLLLOCK,tipd_PLLLOCK);
      VitalWireDelay (RECAL_ipd,RECAL,tipd_RECAL);
      VitalWireDelay (SELFREFRESHENTER_ipd,SELFREFRESHENTER,tipd_SELFREFRESHENTER);
      VitalWireDelay (SYSRST_ipd,SYSRST,tipd_SYSRST);
      VitalWireDelay (UDQSIOIN_ipd,UDQSIOIN,tipd_UDQSIOIN);
      VitalWireDelay (UDQSIOIP_ipd,UDQSIOIP,tipd_UDQSIOIP);
      VitalWireDelay (UIADD_ipd,UIADD,tipd_UIADD);
      VitalWireDelay (UIBROADCAST_ipd,UIBROADCAST,tipd_UIBROADCAST);
      VitalWireDelay (UICLK_ipd,UICLK,tipd_UICLK);
      VitalWireDelay (UICMDEN_ipd,UICMDEN,tipd_UICMDEN);
      VitalWireDelay (UICMDIN_ipd,UICMDIN,tipd_UICMDIN);
      VitalWireDelay (UICMD_ipd,UICMD,tipd_UICMD);
      VitalWireDelay (UICS_ipd,UICS,tipd_UICS);
      VitalWireDelay (UIDONECAL_ipd,UIDONECAL,tipd_UIDONECAL);
      VitalWireDelay (UIDQLOWERDEC_ipd,UIDQLOWERDEC,tipd_UIDQLOWERDEC);
      VitalWireDelay (UIDQLOWERINC_ipd,UIDQLOWERINC,tipd_UIDQLOWERINC);
      VitalWireDelay (UIDQUPPERDEC_ipd,UIDQUPPERDEC,tipd_UIDQUPPERDEC);
      VitalWireDelay (UIDQUPPERINC_ipd,UIDQUPPERINC,tipd_UIDQUPPERINC);
      VitalWireDelay (UIDRPUPDATE_ipd,UIDRPUPDATE,tipd_UIDRPUPDATE);
      VitalWireDelay (UILDQSDEC_ipd,UILDQSDEC,tipd_UILDQSDEC);
      VitalWireDelay (UILDQSINC_ipd,UILDQSINC,tipd_UILDQSINC);
      VitalWireDelay (UIREAD_ipd,UIREAD,tipd_UIREAD);
      VitalWireDelay (UISDI_ipd,UISDI,tipd_UISDI);
      VitalWireDelay (UIUDQSDEC_ipd,UIUDQSDEC,tipd_UIUDQSDEC);
      VitalWireDelay (UIUDQSINC_ipd,UIUDQSINC,tipd_UIUDQSINC);
    end block;
    
    SignalDelay : block
    begin
      P0CMDBA_P0CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P0CMDBA_P0CMDCLK_dly(i),P0CMDBA_ipd(i),tisd_P0CMDBA_P0CMDCLK(i));
      end generate P0CMDBA_P0CMDCLK_DELAY;
      P0CMDBL_P0CMDCLK_DELAY : for i in 5 downto 0 generate
        VitalSignalDelay (P0CMDBL_P0CMDCLK_dly(i),P0CMDBL_ipd(i),tisd_P0CMDBL_P0CMDCLK(i));
      end generate P0CMDBL_P0CMDCLK_DELAY;
      P0CMDCA_P0CMDCLK_DELAY : for i in 11 downto 0 generate
        VitalSignalDelay (P0CMDCA_P0CMDCLK_dly(i),P0CMDCA_ipd(i),tisd_P0CMDCA_P0CMDCLK(i));
      end generate P0CMDCA_P0CMDCLK_DELAY;
      P0CMDINSTR_P0CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P0CMDINSTR_P0CMDCLK_dly(i),P0CMDINSTR_ipd(i),tisd_P0CMDINSTR_P0CMDCLK(i));
      end generate P0CMDINSTR_P0CMDCLK_DELAY;
      P0CMDRA_P0CMDCLK_DELAY : for i in 14 downto 0 generate
        VitalSignalDelay (P0CMDRA_P0CMDCLK_dly(i),P0CMDRA_ipd(i),tisd_P0CMDRA_P0CMDCLK(i));
      end generate P0CMDRA_P0CMDCLK_DELAY;
      P0RWRMASK_P0WRCLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (P0RWRMASK_P0WRCLK_dly(i),P0RWRMASK_ipd(i),tisd_P0RWRMASK_P0WRCLK(i));
      end generate P0RWRMASK_P0WRCLK_DELAY;
      P0WRDATA_P0WRCLK_DELAY : for i in 31 downto 0 generate
        VitalSignalDelay (P0WRDATA_P0WRCLK_dly(i),P0WRDATA_ipd(i),tisd_P0WRDATA_P0WRCLK(i));
      end generate P0WRDATA_P0WRCLK_DELAY;
      P1CMDBA_P1CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P1CMDBA_P1CMDCLK_dly(i),P1CMDBA_ipd(i),tisd_P1CMDBA_P1CMDCLK(i));
      end generate P1CMDBA_P1CMDCLK_DELAY;
      P1CMDBL_P1CMDCLK_DELAY : for i in 5 downto 0 generate
        VitalSignalDelay (P1CMDBL_P1CMDCLK_dly(i),P1CMDBL_ipd(i),tisd_P1CMDBL_P1CMDCLK(i));
      end generate P1CMDBL_P1CMDCLK_DELAY;
      P1CMDCA_P1CMDCLK_DELAY : for i in 11 downto 0 generate
        VitalSignalDelay (P1CMDCA_P1CMDCLK_dly(i),P1CMDCA_ipd(i),tisd_P1CMDCA_P1CMDCLK(i));
      end generate P1CMDCA_P1CMDCLK_DELAY;
      P1CMDINSTR_P1CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P1CMDINSTR_P1CMDCLK_dly(i),P1CMDINSTR_ipd(i),tisd_P1CMDINSTR_P1CMDCLK(i));
      end generate P1CMDINSTR_P1CMDCLK_DELAY;
      P1CMDRA_P1CMDCLK_DELAY : for i in 14 downto 0 generate
        VitalSignalDelay (P1CMDRA_P1CMDCLK_dly(i),P1CMDRA_ipd(i),tisd_P1CMDRA_P1CMDCLK(i));
      end generate P1CMDRA_P1CMDCLK_DELAY;
      P1RWRMASK_P1WRCLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (P1RWRMASK_P1WRCLK_dly(i),P1RWRMASK_ipd(i),tisd_P1RWRMASK_P1WRCLK(i));
      end generate P1RWRMASK_P1WRCLK_DELAY;
      P1WRDATA_P1WRCLK_DELAY : for i in 31 downto 0 generate
        VitalSignalDelay (P1WRDATA_P1WRCLK_dly(i),P1WRDATA_ipd(i),tisd_P1WRDATA_P1WRCLK(i));
      end generate P1WRDATA_P1WRCLK_DELAY;
      P2CMDBA_P2CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P2CMDBA_P2CMDCLK_dly(i),P2CMDBA_ipd(i),tisd_P2CMDBA_P2CMDCLK(i));
      end generate P2CMDBA_P2CMDCLK_DELAY;
      P2CMDBL_P2CMDCLK_DELAY : for i in 5 downto 0 generate
        VitalSignalDelay (P2CMDBL_P2CMDCLK_dly(i),P2CMDBL_ipd(i),tisd_P2CMDBL_P2CMDCLK(i));
      end generate P2CMDBL_P2CMDCLK_DELAY;
      P2CMDCA_P2CMDCLK_DELAY : for i in 11 downto 0 generate
        VitalSignalDelay (P2CMDCA_P2CMDCLK_dly(i),P2CMDCA_ipd(i),tisd_P2CMDCA_P2CMDCLK(i));
      end generate P2CMDCA_P2CMDCLK_DELAY;
      P2CMDINSTR_P2CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P2CMDINSTR_P2CMDCLK_dly(i),P2CMDINSTR_ipd(i),tisd_P2CMDINSTR_P2CMDCLK(i));
      end generate P2CMDINSTR_P2CMDCLK_DELAY;
      P2CMDRA_P2CMDCLK_DELAY : for i in 14 downto 0 generate
        VitalSignalDelay (P2CMDRA_P2CMDCLK_dly(i),P2CMDRA_ipd(i),tisd_P2CMDRA_P2CMDCLK(i));
      end generate P2CMDRA_P2CMDCLK_DELAY;
      P2WRDATA_P2CLK_DELAY : for i in 31 downto 0 generate
        VitalSignalDelay (P2WRDATA_P2CLK_dly(i),P2WRDATA_ipd(i),tisd_P2WRDATA_P2CLK(i));
      end generate P2WRDATA_P2CLK_DELAY;
      P2WRMASK_P2CLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (P2WRMASK_P2CLK_dly(i),P2WRMASK_ipd(i),tisd_P2WRMASK_P2CLK(i));
      end generate P2WRMASK_P2CLK_DELAY;
      P3CMDBA_P3CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P3CMDBA_P3CMDCLK_dly(i),P3CMDBA_ipd(i),tisd_P3CMDBA_P3CMDCLK(i));
      end generate P3CMDBA_P3CMDCLK_DELAY;
      P3CMDBL_P3CMDCLK_DELAY : for i in 5 downto 0 generate
        VitalSignalDelay (P3CMDBL_P3CMDCLK_dly(i),P3CMDBL_ipd(i),tisd_P3CMDBL_P3CMDCLK(i));
      end generate P3CMDBL_P3CMDCLK_DELAY;
      P3CMDCA_P3CMDCLK_DELAY : for i in 11 downto 0 generate
        VitalSignalDelay (P3CMDCA_P3CMDCLK_dly(i),P3CMDCA_ipd(i),tisd_P3CMDCA_P3CMDCLK(i));
      end generate P3CMDCA_P3CMDCLK_DELAY;
      P3CMDINSTR_P3CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P3CMDINSTR_P3CMDCLK_dly(i),P3CMDINSTR_ipd(i),tisd_P3CMDINSTR_P3CMDCLK(i));
      end generate P3CMDINSTR_P3CMDCLK_DELAY;
      P3CMDRA_P3CMDCLK_DELAY : for i in 14 downto 0 generate
        VitalSignalDelay (P3CMDRA_P3CMDCLK_dly(i),P3CMDRA_ipd(i),tisd_P3CMDRA_P3CMDCLK(i));
      end generate P3CMDRA_P3CMDCLK_DELAY;
      P3WRDATA_P3CLK_DELAY : for i in 31 downto 0 generate
        VitalSignalDelay (P3WRDATA_P3CLK_dly(i),P3WRDATA_ipd(i),tisd_P3WRDATA_P3CLK(i));
      end generate P3WRDATA_P3CLK_DELAY;
      P3WRMASK_P3CLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (P3WRMASK_P3CLK_dly(i),P3WRMASK_ipd(i),tisd_P3WRMASK_P3CLK(i));
      end generate P3WRMASK_P3CLK_DELAY;
      P4CMDBA_P4CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P4CMDBA_P4CMDCLK_dly(i),P4CMDBA_ipd(i),tisd_P4CMDBA_P4CMDCLK(i));
      end generate P4CMDBA_P4CMDCLK_DELAY;
      P4CMDBL_P4CMDCLK_DELAY : for i in 5 downto 0 generate
        VitalSignalDelay (P4CMDBL_P4CMDCLK_dly(i),P4CMDBL_ipd(i),tisd_P4CMDBL_P4CMDCLK(i));
      end generate P4CMDBL_P4CMDCLK_DELAY;
      P4CMDCA_P4CMDCLK_DELAY : for i in 11 downto 0 generate
        VitalSignalDelay (P4CMDCA_P4CMDCLK_dly(i),P4CMDCA_ipd(i),tisd_P4CMDCA_P4CMDCLK(i));
      end generate P4CMDCA_P4CMDCLK_DELAY;
      P4CMDINSTR_P4CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P4CMDINSTR_P4CMDCLK_dly(i),P4CMDINSTR_ipd(i),tisd_P4CMDINSTR_P4CMDCLK(i));
      end generate P4CMDINSTR_P4CMDCLK_DELAY;
      P4CMDRA_P4CMDCLK_DELAY : for i in 14 downto 0 generate
        VitalSignalDelay (P4CMDRA_P4CMDCLK_dly(i),P4CMDRA_ipd(i),tisd_P4CMDRA_P4CMDCLK(i));
      end generate P4CMDRA_P4CMDCLK_DELAY;
      P4WRDATA_P4CLK_DELAY : for i in 31 downto 0 generate
        VitalSignalDelay (P4WRDATA_P4CLK_dly(i),P4WRDATA_ipd(i),tisd_P4WRDATA_P4CLK(i));
      end generate P4WRDATA_P4CLK_DELAY;
      P4WRMASK_P4CLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (P4WRMASK_P4CLK_dly(i),P4WRMASK_ipd(i),tisd_P4WRMASK_P4CLK(i));
      end generate P4WRMASK_P4CLK_DELAY;
      P5CMDBA_P5CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P5CMDBA_P5CMDCLK_dly(i),P5CMDBA_ipd(i),tisd_P5CMDBA_P5CMDCLK(i));
      end generate P5CMDBA_P5CMDCLK_DELAY;
      P5CMDBL_P5CMDCLK_DELAY : for i in 5 downto 0 generate
        VitalSignalDelay (P5CMDBL_P5CMDCLK_dly(i),P5CMDBL_ipd(i),tisd_P5CMDBL_P5CMDCLK(i));
      end generate P5CMDBL_P5CMDCLK_DELAY;
      P5CMDCA_P5CMDCLK_DELAY : for i in 11 downto 0 generate
        VitalSignalDelay (P5CMDCA_P5CMDCLK_dly(i),P5CMDCA_ipd(i),tisd_P5CMDCA_P5CMDCLK(i));
      end generate P5CMDCA_P5CMDCLK_DELAY;
      P5CMDINSTR_P5CMDCLK_DELAY : for i in 2 downto 0 generate
        VitalSignalDelay (P5CMDINSTR_P5CMDCLK_dly(i),P5CMDINSTR_ipd(i),tisd_P5CMDINSTR_P5CMDCLK(i));
      end generate P5CMDINSTR_P5CMDCLK_DELAY;
      P5CMDRA_P5CMDCLK_DELAY : for i in 14 downto 0 generate
        VitalSignalDelay (P5CMDRA_P5CMDCLK_dly(i),P5CMDRA_ipd(i),tisd_P5CMDRA_P5CMDCLK(i));
      end generate P5CMDRA_P5CMDCLK_DELAY;
      P5WRDATA_P5CLK_DELAY : for i in 31 downto 0 generate
        VitalSignalDelay (P5WRDATA_P5CLK_dly(i),P5WRDATA_ipd(i),tisd_P5WRDATA_P5CLK(i));
      end generate P5WRDATA_P5CLK_DELAY;
      P5WRMASK_P5CLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (P5WRMASK_P5CLK_dly(i),P5WRMASK_ipd(i),tisd_P5WRMASK_P5CLK(i));
      end generate P5WRMASK_P5CLK_DELAY;
      PLLCE_PLLCLK_DELAY_0 : for i in 1 downto 0 generate
        VitalSignalDelay (PLLCE_PLLCLK_dly(i),PLLCE_ipd(0),tisd_PLLCE_PLLCLK(i));
      end generate PLLCE_PLLCLK_DELAY_0;
      PLLCE_PLLCLK_DELAY_1 : for i in 3 downto 2 generate
        VitalSignalDelay (PLLCE_PLLCLK_dly(i),PLLCE_ipd(1),tisd_PLLCE_PLLCLK(i));
      end generate PLLCE_PLLCLK_DELAY_1;
      PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (PLLCLK_dly(i),PLLCLK_ipd(i),ticd_PLLCLK(i));
      end generate PLLCLK_DELAY;
      UIADDR_UICLK_DELAY : for i in 4 downto 0 generate
        VitalSignalDelay (UIADDR_UICLK_dly(i),UIADDR_ipd(i),tisd_UIADDR_UICLK(i));
      end generate UIADDR_UICLK_DELAY;
      UIDQCOUNT_UICLK_DELAY : for i in 3 downto 0 generate
        VitalSignalDelay (UIDQCOUNT_UICLK_dly(i),UIDQCOUNT_ipd(i),tisd_UIDQCOUNT_UICLK(i));
      end generate UIDQCOUNT_UICLK_DELAY;
      VitalSignalDelay (IOIDRPSDI_UICLK_dly,IOIDRPSDI_ipd,tisd_IOIDRPSDI_UICLK);
      P0ARBEN_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (P0ARBEN_PLLCLK_dly(i),P0ARBEN_ipd,tisd_P0ARBEN_PLLCLK(i));
      end generate P0ARBEN_PLLCLK_DELAY;
      VitalSignalDelay (P0CMDEN_P0CMDCLK_dly,P0CMDEN_ipd,tisd_P0CMDEN_P0CMDCLK);
      VitalSignalDelay (P0RDEN_P0RDCLK_dly,P0RDEN_ipd,tisd_P0RDEN_P0RDCLK);
      VitalSignalDelay (P0WREN_P0WRCLK_dly,P0WREN_ipd,tisd_P0WREN_P0WRCLK);
      P1ARBEN_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (P1ARBEN_PLLCLK_dly(i),P1ARBEN_ipd,tisd_P1ARBEN_PLLCLK(i));
      end generate P1ARBEN_PLLCLK_DELAY;
      VitalSignalDelay (P1CMDEN_P1CMDCLK_dly,P1CMDEN_ipd,tisd_P1CMDEN_P1CMDCLK);
      VitalSignalDelay (P1RDEN_P1RDCLK_dly,P1RDEN_ipd,tisd_P1RDEN_P1RDCLK);
      VitalSignalDelay (P1WREN_P1WRCLK_dly,P1WREN_ipd,tisd_P1WREN_P1WRCLK);
      P2ARBEN_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (P2ARBEN_PLLCLK_dly(i),P2ARBEN_ipd,tisd_P2ARBEN_PLLCLK(i));
      end generate P2ARBEN_PLLCLK_DELAY;
      VitalSignalDelay (P2CMDEN_P2CMDCLK_dly,P2CMDEN_ipd,tisd_P2CMDEN_P2CMDCLK);
      VitalSignalDelay (P2EN_P2CLK_dly,P2EN_ipd,tisd_P2EN_P2CLK);
      P3ARBEN_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (P3ARBEN_PLLCLK_dly(i),P3ARBEN_ipd,tisd_P3ARBEN_PLLCLK(i));
      end generate P3ARBEN_PLLCLK_DELAY;
      VitalSignalDelay (P3CMDEN_P3CMDCLK_dly,P3CMDEN_ipd,tisd_P3CMDEN_P3CMDCLK);
      VitalSignalDelay (P3EN_P3CLK_dly,P3EN_ipd,tisd_P3EN_P3CLK);
      P4ARBEN_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (P4ARBEN_PLLCLK_dly(i),P4ARBEN_ipd,tisd_P4ARBEN_PLLCLK(i));
      end generate P4ARBEN_PLLCLK_DELAY;
      VitalSignalDelay (P4CMDEN_P4CMDCLK_dly,P4CMDEN_ipd,tisd_P4CMDEN_P4CMDCLK);
      VitalSignalDelay (P4EN_P4CLK_dly,P4EN_ipd,tisd_P4EN_P4CLK);
      P5ARBEN_PLLCLK_DELAY : for i in 1 downto 0 generate
       VitalSignalDelay (P5ARBEN_PLLCLK_dly(i),P5ARBEN_ipd,tisd_P5ARBEN_PLLCLK(i));
      end generate P5ARBEN_PLLCLK_DELAY;
      VitalSignalDelay (P5CMDEN_P5CMDCLK_dly,P5CMDEN_ipd,tisd_P5CMDEN_P5CMDCLK);
      VitalSignalDelay (P5EN_P5CLK_dly,P5EN_ipd,tisd_P5EN_P5CLK);
      PLLLOCK_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (PLLLOCK_PLLCLK_dly(i),PLLLOCK_ipd,tisd_PLLLOCK_PLLCLK(i));
      end generate PLLLOCK_PLLCLK_DELAY;
      RECAL_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (RECAL_PLLCLK_dly(i),RECAL_ipd,tisd_RECAL_PLLCLK(i));
      end generate RECAL_PLLCLK_DELAY;
      SELFREFRESHENTER_PLLCLK_DELAY : for i in 1 downto 0 generate
        VitalSignalDelay (SELFREFRESHENTER_PLLCLK_dly(i),SELFREFRESHENTER_ipd,tisd_SELFREFRESHENTER_PLLCLK(i));
      end generate SELFREFRESHENTER_PLLCLK_DELAY;
      VitalSignalDelay (UIADD_UICLK_dly,UIADD_ipd,tisd_UIADD_UICLK);
      VitalSignalDelay (UIBROADCAST_UICLK_dly,UIBROADCAST_ipd,tisd_UIBROADCAST_UICLK);
      VitalSignalDelay (UICMDEN_UICLK_dly,UICMDEN_ipd,tisd_UICMDEN_UICLK);
      VitalSignalDelay (UICMDIN_UICLK_dly,UICMDIN_ipd,tisd_UICMDIN_UICLK);
      VitalSignalDelay (UICMD_UICLK_dly,UICMD_ipd,tisd_UICMD_UICLK);
      VitalSignalDelay (UICS_UICLK_dly,UICS_ipd,tisd_UICS_UICLK);
      VitalSignalDelay (UIDONECAL_UICLK_dly,UIDONECAL_ipd,tisd_UIDONECAL_UICLK);
      VitalSignalDelay (UIDQLOWERDEC_UICLK_dly,UIDQLOWERDEC_ipd,tisd_UIDQLOWERDEC_UICLK);
      VitalSignalDelay (UIDQLOWERINC_UICLK_dly,UIDQLOWERINC_ipd,tisd_UIDQLOWERINC_UICLK);
      VitalSignalDelay (UIDQUPPERDEC_UICLK_dly,UIDQUPPERDEC_ipd,tisd_UIDQUPPERDEC_UICLK);
      VitalSignalDelay (UIDQUPPERINC_UICLK_dly,UIDQUPPERINC_ipd,tisd_UIDQUPPERINC_UICLK);
      VitalSignalDelay (UIDRPUPDATE_UICLK_dly,UIDRPUPDATE_ipd,tisd_UIDRPUPDATE_UICLK);
      VitalSignalDelay (UILDQSDEC_UICLK_dly,UILDQSDEC_ipd,tisd_UILDQSDEC_UICLK);
      VitalSignalDelay (UILDQSINC_UICLK_dly,UILDQSINC_ipd,tisd_UILDQSINC_UICLK);
      VitalSignalDelay (UIREAD_UICLK_dly,UIREAD_ipd,tisd_UIREAD_UICLK);
      VitalSignalDelay (UISDI_UICLK_dly,UISDI_ipd,tisd_UISDI_UICLK);
      VitalSignalDelay (UIUDQSDEC_UICLK_dly,UIUDQSDEC_ipd,tisd_UIUDQSDEC_UICLK);
      VitalSignalDelay (UIUDQSINC_UICLK_dly,UIUDQSINC_ipd,tisd_UIUDQSINC_UICLK);

      VitalSignalDelay (P0CMDCLK_dly,P0CMDCLK_ipd,ticd_P0CMDCLK);
      VitalSignalDelay (P0RDCLK_dly,P0RDCLK_ipd,ticd_P0RDCLK);
      VitalSignalDelay (P0WRCLK_dly,P0WRCLK_ipd,ticd_P0WRCLK);
      VitalSignalDelay (P1CMDCLK_dly,P1CMDCLK_ipd,ticd_P1CMDCLK);
      VitalSignalDelay (P1RDCLK_dly,P1RDCLK_ipd,ticd_P1RDCLK);
      VitalSignalDelay (P1WRCLK_dly,P1WRCLK_ipd,ticd_P1WRCLK);
      VitalSignalDelay (P2CLK_dly,P2CLK_ipd,ticd_P2CLK);
      VitalSignalDelay (P2CMDCLK_dly,P2CMDCLK_ipd,ticd_P2CMDCLK);
      VitalSignalDelay (P3CLK_dly,P3CLK_ipd,ticd_P3CLK);
      VitalSignalDelay (P3CMDCLK_dly,P3CMDCLK_ipd,ticd_P3CMDCLK);
      VitalSignalDelay (P4CLK_dly,P4CLK_ipd,ticd_P4CLK);
      VitalSignalDelay (P4CMDCLK_dly,P4CMDCLK_ipd,ticd_P4CMDCLK);
      VitalSignalDelay (P5CLK_dly,P5CLK_ipd,ticd_P5CLK);
      VitalSignalDelay (P5CMDCLK_dly,P5CMDCLK_ipd,ticd_P5CMDCLK);
      VitalSignalDelay (UICLK_dly,UICLK_ipd,ticd_UICLK);
    end block;

    SELECTPROC : process(P0ARBEN_PLLCLK_dly, P1ARBEN_PLLCLK_dly, P2ARBEN_PLLCLK_dly, P3ARBEN_PLLCLK_dly, P4ARBEN_PLLCLK_dly, P5ARBEN_PLLCLK_dly, 
                         PLLLOCK_PLLCLK_dly, RECAL_PLLCLK_dly, SELFREFRESHENTER_PLLCLK_dly, PLLCE_PLLCLK_dly)
    begin 
      if(abs(tisd_P0ARBEN_PLLCLK(0))> abs(tisd_P0ARBEN_PLLCLK(1))) then
        P0ARBEN_indelay <= P0ARBEN_PLLCLK_dly(0);
        else
        P0ARBEN_indelay <= P0ARBEN_PLLCLK_dly(1);
      end if;
      if(abs(tisd_P1ARBEN_PLLCLK(0))> abs(tisd_P1ARBEN_PLLCLK(1))) then
        P1ARBEN_indelay <= P1ARBEN_PLLCLK_dly(0);
        else
        P1ARBEN_indelay <= P1ARBEN_PLLCLK_dly(1);
      end if;
      if(abs(tisd_P2ARBEN_PLLCLK(0))> abs(tisd_P2ARBEN_PLLCLK(1))) then
        P2ARBEN_indelay <= P2ARBEN_PLLCLK_dly(0);
        else
        P2ARBEN_indelay <= P2ARBEN_PLLCLK_dly(1);
      end if;
      if(abs(tisd_P3ARBEN_PLLCLK(0))> abs(tisd_P3ARBEN_PLLCLK(1))) then
        P3ARBEN_indelay <= P3ARBEN_PLLCLK_dly(0);
        else
        P3ARBEN_indelay <= P3ARBEN_PLLCLK_dly(1);
      end if;
      if(abs(tisd_P4ARBEN_PLLCLK(0))> abs(tisd_P4ARBEN_PLLCLK(1))) then
        P4ARBEN_indelay <= P4ARBEN_PLLCLK_dly(0);
        else
        P4ARBEN_indelay <= P4ARBEN_PLLCLK_dly(1);
      end if;
      if(abs(tisd_P5ARBEN_PLLCLK(0))> abs(tisd_P5ARBEN_PLLCLK(1))) then
        P5ARBEN_indelay <= P5ARBEN_PLLCLK_dly(0);
        else
        P5ARBEN_indelay <= P5ARBEN_PLLCLK_dly(1);
      end if;
      if(abs(tisd_PLLLOCK_PLLCLK(0))> abs(tisd_PLLLOCK_PLLCLK(1))) then
        PLLLOCK_indelay <= PLLLOCK_PLLCLK_dly(0);
        else
        PLLLOCK_indelay <= PLLLOCK_PLLCLK_dly(1);
      end if;
      if(abs(tisd_RECAL_PLLCLK(0))> abs(tisd_RECAL_PLLCLK(1))) then
        RECAL_indelay <= RECAL_PLLCLK_dly(0);
        else
        RECAL_indelay <= RECAL_PLLCLK_dly(1);
      end if;
      if(abs(tisd_SELFREFRESHENTER_PLLCLK(0))> abs(tisd_SELFREFRESHENTER_PLLCLK(1))) then
        SELFREFRESHENTER_indelay <= SELFREFRESHENTER_PLLCLK_dly(0);
        else
        SELFREFRESHENTER_indelay <= SELFREFRESHENTER_PLLCLK_dly(1);
      end if;
      if(abs(tisd_PLLCE_PLLCLK(0)) > tisd_PLLCE_PLLCLK(1)) then
        PLLCE_indelay(0) <= PLLCE_PLLCLK_dly(0);
      else
        PLLCE_indelay(0) <= PLLCE_PLLCLK_dly(1);
      end if;
      if(abs(tisd_PLLCE_PLLCLK(2)) > tisd_PLLCE_PLLCLK(3)) then
        PLLCE_indelay(1) <= PLLCE_PLLCLK_dly(2);
      else
        PLLCE_indelay(1) <= PLLCE_PLLCLK_dly(3);
      end if;
    end process;

    --Input ports sensitive to single clock
    IOIDRPSDI_indelay <= IOIDRPSDI_UICLK_dly;
    P0CMDBA_indelay <= P0CMDBA_P0CMDCLK_dly;
    P0CMDBL_indelay <= P0CMDBL_P0CMDCLK_dly;
    P0CMDCA_indelay <= P0CMDCA_P0CMDCLK_dly;
    P0CMDEN_indelay <= P0CMDEN_P0CMDCLK_dly;
    P0CMDINSTR_indelay <= P0CMDINSTR_P0CMDCLK_dly;
    P0CMDRA_indelay <= P0CMDRA_P0CMDCLK_dly;
    P0RDEN_indelay <= P0RDEN_P0RDCLK_dly;
    P0RWRMASK_indelay <= P0RWRMASK_P0WRCLK_dly;
    P0WRDATA_indelay <= P0WRDATA_P0WRCLK_dly;
    P0WREN_indelay <= P0WREN_P0WRCLK_dly;
    P1CMDBA_indelay <= P1CMDBA_P1CMDCLK_dly;
    P1CMDBL_indelay <= P1CMDBL_P1CMDCLK_dly;
    P1CMDCA_indelay <= P1CMDCA_P1CMDCLK_dly;
    P1CMDEN_indelay <= P1CMDEN_P1CMDCLK_dly;
    P1CMDINSTR_indelay <= P1CMDINSTR_P1CMDCLK_dly;
    P1CMDRA_indelay <= P1CMDRA_P1CMDCLK_dly;
    P1RDEN_indelay <= P1RDEN_P1RDCLK_dly;
    P1RWRMASK_indelay <= P1RWRMASK_P1WRCLK_dly;
    P1WRDATA_indelay <= P1WRDATA_P1WRCLK_dly;
    P1WREN_indelay <= P1WREN_P1WRCLK_dly;
    P2CMDBA_indelay <= P2CMDBA_P2CMDCLK_dly;
    P2CMDBL_indelay <= P2CMDBL_P2CMDCLK_dly;
    P2CMDCA_indelay <= P2CMDCA_P2CMDCLK_dly;
    P2CMDEN_indelay <= P2CMDEN_P2CMDCLK_dly;
    P2CMDINSTR_indelay <= P2CMDINSTR_P2CMDCLK_dly;
    P2CMDRA_indelay <= P2CMDRA_P2CMDCLK_dly;
    P2EN_indelay <= P2EN_P2CLK_dly;
    P2WRDATA_indelay <= P2WRDATA_P2CLK_dly;
    P2WRMASK_indelay <= P2WRMASK_P2CLK_dly;
    P3CMDBA_indelay <= P3CMDBA_P3CMDCLK_dly;
    P3CMDBL_indelay <= P3CMDBL_P3CMDCLK_dly;
    P3CMDCA_indelay <= P3CMDCA_P3CMDCLK_dly;
    P3CMDEN_indelay <= P3CMDEN_P3CMDCLK_dly;
    P3CMDINSTR_indelay <= P3CMDINSTR_P3CMDCLK_dly;
    P3CMDRA_indelay <= P3CMDRA_P3CMDCLK_dly;
    P3EN_indelay <= P3EN_P3CLK_dly;
    P3WRDATA_indelay <= P3WRDATA_P3CLK_dly;
    P3WRMASK_indelay <= P3WRMASK_P3CLK_dly;
    P4CMDBA_indelay <= P4CMDBA_P4CMDCLK_dly;
    P4CMDBL_indelay <= P4CMDBL_P4CMDCLK_dly;
    P4CMDCA_indelay <= P4CMDCA_P4CMDCLK_dly;
    P4CMDEN_indelay <= P4CMDEN_P4CMDCLK_dly;
    P4CMDINSTR_indelay <= P4CMDINSTR_P4CMDCLK_dly;
    P4CMDRA_indelay <= P4CMDRA_P4CMDCLK_dly;
    P4EN_indelay <= P4EN_P4CLK_dly;
    P4WRDATA_indelay <= P4WRDATA_P4CLK_dly;
    P4WRMASK_indelay <= P4WRMASK_P4CLK_dly;
    P5CMDBA_indelay <= P5CMDBA_P5CMDCLK_dly;
    P5CMDBL_indelay <= P5CMDBL_P5CMDCLK_dly;
    P5CMDCA_indelay <= P5CMDCA_P5CMDCLK_dly;
    P5CMDEN_indelay <= P5CMDEN_P5CMDCLK_dly;
    P5CMDINSTR_indelay <= P5CMDINSTR_P5CMDCLK_dly;
    P5CMDRA_indelay <= P5CMDRA_P5CMDCLK_dly;
    P5EN_indelay <= P5EN_P5CLK_dly;
    P5WRDATA_indelay <= P5WRDATA_P5CLK_dly;
    P5WRMASK_indelay <= P5WRMASK_P5CLK_dly;
    UIADDR_indelay <= UIADDR_UICLK_dly;
    UIADD_indelay <= UIADD_UICLK_dly;
    UIBROADCAST_indelay <= UIBROADCAST_UICLK_dly;
    UICMDEN_indelay <= UICMDEN_UICLK_dly;
    UICMDIN_indelay <= UICMDIN_UICLK_dly;
    UICMD_indelay <= UICMD_UICLK_dly;
    UICS_indelay <= UICS_UICLK_dly;
    UIDONECAL_indelay <= UIDONECAL_UICLK_dly;
    UIDQCOUNT_indelay <= UIDQCOUNT_UICLK_dly;
    UIDQLOWERDEC_indelay <= UIDQLOWERDEC_UICLK_dly;
    UIDQLOWERINC_indelay <= UIDQLOWERINC_UICLK_dly;
    UIDQUPPERDEC_indelay <= UIDQUPPERDEC_UICLK_dly;
    UIDQUPPERINC_indelay <= UIDQUPPERINC_UICLK_dly;
    UIDRPUPDATE_indelay <= UIDRPUPDATE_UICLK_dly;
    UILDQSDEC_indelay <= UILDQSDEC_UICLK_dly;
    UILDQSINC_indelay <= UILDQSINC_UICLK_dly;
    UIREAD_indelay <= UIREAD_UICLK_dly;
    UISDI_indelay <= UISDI_UICLK_dly;
    UIUDQSDEC_indelay <= UIUDQSDEC_UICLK_dly;
    UIUDQSINC_indelay <= UIUDQSINC_UICLK_dly;
    
    DQI_indelay <= DQI_ipd;
    DQSIOIN_indelay <= DQSIOIN_ipd;
    DQSIOIP_indelay <= DQSIOIP_ipd;
    SYSRST_indelay <= SYSRST_ipd;
    UDQSIOIN_indelay <= UDQSIOIN_ipd;
    UDQSIOIP_indelay <= UDQSIOIP_ipd;
    
    P0CMDCLK_indelay <= P0CMDCLK_dly;
    P0RDCLK_indelay <= P0RDCLK_dly;
    P0WRCLK_indelay <= P0WRCLK_dly;
    P1CMDCLK_indelay <= P1CMDCLK_dly;
    P1RDCLK_indelay <= P1RDCLK_dly;
    P1WRCLK_indelay <= P1WRCLK_dly;
    P2CLK_indelay <= P2CLK_dly;
    P2CMDCLK_indelay <= P2CMDCLK_dly;
    P3CLK_indelay <= P3CLK_dly;
    P3CMDCLK_indelay <= P3CMDCLK_dly;
    P4CLK_indelay <= P4CLK_dly;
    P4CMDCLK_indelay <= P4CMDCLK_dly;
    P5CLK_indelay <= P5CLK_dly;
    P5CMDCLK_indelay <= P5CMDCLK_dly;
    PLLCLK_indelay <= PLLCLK_dly;
    UICLK_indelay <= UICLK_dly;
    
    ADDR_out <= ADDR_outdelay after OUT_DELAY;
    BA_out <= BA_outdelay after OUT_DELAY;
    CAS_out <= CAS_outdelay after OUT_DELAY;
    CKE_out <= CKE_outdelay after OUT_DELAY;
    DQIOWEN0_out <= DQIOWEN0_outdelay after OUT_DELAY;
    DQON_out <= DQON_outdelay after OUT_DELAY;
    DQOP_out <= DQOP_outdelay after OUT_DELAY;
    DQSIOWEN90N_out <= DQSIOWEN90N_outdelay after OUT_DELAY;
    DQSIOWEN90P_out <= DQSIOWEN90P_outdelay after OUT_DELAY;
    IOIDRPADDR_out <= IOIDRPADDR_outdelay after OUT_DELAY;
    IOIDRPADD_out <= IOIDRPADD_outdelay after OUT_DELAY;
    IOIDRPBROADCAST_out <= IOIDRPBROADCAST_outdelay after OUT_DELAY;
    IOIDRPCLK_out <= IOIDRPCLK_outdelay after 0 ps;
    IOIDRPCS_out <= IOIDRPCS_outdelay after OUT_DELAY;
    IOIDRPSDO_out <= IOIDRPSDO_outdelay after OUT_DELAY;
    IOIDRPTRAIN_out <= IOIDRPTRAIN_outdelay after OUT_DELAY;
    IOIDRPUPDATE_out <= IOIDRPUPDATE_outdelay after OUT_DELAY;
    LDMN_out <= LDMN_outdelay after OUT_DELAY;
    LDMP_out <= LDMP_outdelay after OUT_DELAY;
    ODT_out <= ODT_outdelay after OUT_DELAY;
    P0CMDEMPTY_out <= P0CMDEMPTY_outdelay after OUT_DELAY;
    P0CMDFULL_out <= P0CMDFULL_outdelay after OUT_DELAY;
    P0RDCOUNT_out <= P0RDCOUNT_outdelay after OUT_DELAY;
    P0RDDATA_out <= P0RDDATA_outdelay after OUT_DELAY;
    P0RDEMPTY_out <= P0RDEMPTY_outdelay after OUT_DELAY;
    P0RDERROR_out <= P0RDERROR_outdelay after OUT_DELAY;
    P0RDFULL_out <= P0RDFULL_outdelay after OUT_DELAY;
    P0RDOVERFLOW_out <= P0RDOVERFLOW_outdelay after OUT_DELAY;
    P0WRCOUNT_out <= P0WRCOUNT_outdelay after OUT_DELAY;
    P0WREMPTY_out <= P0WREMPTY_outdelay after OUT_DELAY;
    P0WRERROR_out <= P0WRERROR_outdelay after OUT_DELAY;
    P0WRFULL_out <= P0WRFULL_outdelay after OUT_DELAY;
    P0WRUNDERRUN_out <= P0WRUNDERRUN_outdelay after OUT_DELAY;
    P1CMDEMPTY_out <= P1CMDEMPTY_outdelay after OUT_DELAY;
    P1CMDFULL_out <= P1CMDFULL_outdelay after OUT_DELAY;
    P1RDCOUNT_out <= P1RDCOUNT_outdelay after OUT_DELAY;
    P1RDDATA_out <= P1RDDATA_outdelay after OUT_DELAY;
    P1RDEMPTY_out <= P1RDEMPTY_outdelay after OUT_DELAY;
    P1RDERROR_out <= P1RDERROR_outdelay after OUT_DELAY;
    P1RDFULL_out <= P1RDFULL_outdelay after OUT_DELAY;
    P1RDOVERFLOW_out <= P1RDOVERFLOW_outdelay after OUT_DELAY;
    P1WRCOUNT_out <= P1WRCOUNT_outdelay after OUT_DELAY;
    P1WREMPTY_out <= P1WREMPTY_outdelay after OUT_DELAY;
    P1WRERROR_out <= P1WRERROR_outdelay after OUT_DELAY;
    P1WRFULL_out <= P1WRFULL_outdelay after OUT_DELAY;
    P1WRUNDERRUN_out <= P1WRUNDERRUN_outdelay after OUT_DELAY;
    P2CMDEMPTY_out <= P2CMDEMPTY_outdelay after OUT_DELAY;
    P2CMDFULL_out <= P2CMDFULL_outdelay after OUT_DELAY;
    P2COUNT_out <= P2COUNT_outdelay after OUT_DELAY;
    P2EMPTY_out <= P2EMPTY_outdelay after OUT_DELAY;
    P2ERROR_out <= P2ERROR_outdelay after OUT_DELAY;
    P2FULL_out <= P2FULL_outdelay after OUT_DELAY;
    P2RDDATA_out <= P2RDDATA_outdelay after OUT_DELAY;
    P2RDOVERFLOW_out <= P2RDOVERFLOW_outdelay after OUT_DELAY;
    P2WRUNDERRUN_out <= P2WRUNDERRUN_outdelay after OUT_DELAY;
    P3CMDEMPTY_out <= P3CMDEMPTY_outdelay after OUT_DELAY;
    P3CMDFULL_out <= P3CMDFULL_outdelay after OUT_DELAY;
    P3COUNT_out <= P3COUNT_outdelay after OUT_DELAY;
    P3EMPTY_out <= P3EMPTY_outdelay after OUT_DELAY;
    P3ERROR_out <= P3ERROR_outdelay after OUT_DELAY;
    P3FULL_out <= P3FULL_outdelay after OUT_DELAY;
    P3RDDATA_out <= P3RDDATA_outdelay after OUT_DELAY;
    P3RDOVERFLOW_out <= P3RDOVERFLOW_outdelay after OUT_DELAY;
    P3WRUNDERRUN_out <= P3WRUNDERRUN_outdelay after OUT_DELAY;
    P4CMDEMPTY_out <= P4CMDEMPTY_outdelay after OUT_DELAY;
    P4CMDFULL_out <= P4CMDFULL_outdelay after OUT_DELAY;
    P4COUNT_out <= P4COUNT_outdelay after OUT_DELAY;
    P4EMPTY_out <= P4EMPTY_outdelay after OUT_DELAY;
    P4ERROR_out <= P4ERROR_outdelay after OUT_DELAY;
    P4FULL_out <= P4FULL_outdelay after OUT_DELAY;
    P4RDDATA_out <= P4RDDATA_outdelay after OUT_DELAY;
    P4RDOVERFLOW_out <= P4RDOVERFLOW_outdelay after OUT_DELAY;
    P4WRUNDERRUN_out <= P4WRUNDERRUN_outdelay after OUT_DELAY;
    P5CMDEMPTY_out <= P5CMDEMPTY_outdelay after OUT_DELAY;
    P5CMDFULL_out <= P5CMDFULL_outdelay after OUT_DELAY;
    P5COUNT_out <= P5COUNT_outdelay after OUT_DELAY;
    P5EMPTY_out <= P5EMPTY_outdelay after OUT_DELAY;
    P5ERROR_out <= P5ERROR_outdelay after OUT_DELAY;
    P5FULL_out <= P5FULL_outdelay after OUT_DELAY;
    P5RDDATA_out <= P5RDDATA_outdelay after OUT_DELAY;
    P5RDOVERFLOW_out <= P5RDOVERFLOW_outdelay after OUT_DELAY;
    P5WRUNDERRUN_out <= P5WRUNDERRUN_outdelay after OUT_DELAY;
    RAS_out <= RAS_outdelay after OUT_DELAY;
    RST_out <= RST_outdelay after OUT_DELAY;
    SELFREFRESHMODE_out <= SELFREFRESHMODE_outdelay after OUT_DELAY;
    STATUS_out <= STATUS_outdelay after OUT_DELAY;
    UDMN_out <= UDMN_outdelay after OUT_DELAY;
    UDMP_out <= UDMP_outdelay after OUT_DELAY;
    UOCALSTART_out <= UOCALSTART_outdelay after OUT_DELAY;
    UOCMDREADYIN_out <= UOCMDREADYIN_outdelay after OUT_DELAY;
    UODATAVALID_out <= UODATAVALID_outdelay after OUT_DELAY;
    UODATA_out <= UODATA_outdelay after OUT_DELAY;
    UODONECAL_out <= UODONECAL_outdelay after OUT_DELAY;
    UOREFRSHFLAG_out <= UOREFRSHFLAG_outdelay after OUT_DELAY;
    UOSDO_out <= UOSDO_outdelay after OUT_DELAY;
    WE_out <= WE_outdelay after OUT_DELAY;
    
    DQSIOIN_indly <= DQSIOIN_indelay after INCLK_DELAY;
    DQSIOIP_indly <= DQSIOIP_indelay after INCLK_DELAY;
    P0CMDCLK_indly <= P0CMDCLK_indelay after INCLK_DELAY;
    P0RDCLK_indly <= P0RDCLK_indelay after INCLK_DELAY;
    P0WRCLK_indly <= P0WRCLK_indelay after INCLK_DELAY;
    P1CMDCLK_indly <= P1CMDCLK_indelay after INCLK_DELAY;
    P1RDCLK_indly <= P1RDCLK_indelay after INCLK_DELAY;
    P1WRCLK_indly <= P1WRCLK_indelay after INCLK_DELAY;
    P2CLK_indly <= P2CLK_indelay after INCLK_DELAY;
    P2CMDCLK_indly <= P2CMDCLK_indelay after INCLK_DELAY;
    P3CLK_indly <= P3CLK_indelay after INCLK_DELAY;
    P3CMDCLK_indly <= P3CMDCLK_indelay after INCLK_DELAY;
    P4CLK_indly <= P4CLK_indelay after INCLK_DELAY;
    P4CMDCLK_indly <= P4CMDCLK_indelay after INCLK_DELAY;
    P5CLK_indly <= P5CLK_indelay after INCLK_DELAY;
    P5CMDCLK_indly <= P5CMDCLK_indelay after INCLK_DELAY;
    PLLCLK_indly <= PLLCLK_indelay after INCLK_DELAY;
    UDQSIOIN_indly <= UDQSIOIN_indelay after INCLK_DELAY;
    UDQSIOIP_indly <= UDQSIOIP_indelay after INCLK_DELAY;
    UICLK_indly <= UICLK_indelay after INCLK_DELAY;
    
    DQI_indly <= DQI_indelay after IN_DELAY;
    IOIDRPSDI_indly <= IOIDRPSDI_indelay after IN_DELAY;
    P0ARBEN_indly <= P0ARBEN_indelay after IN_DELAY;
    P0CMDBA_indly <= P0CMDBA_indelay after IN_DELAY;
    P0CMDBL_indly <= P0CMDBL_indelay after IN_DELAY;
    P0CMDCA_indly <= P0CMDCA_indelay after IN_DELAY;
    P0CMDEN_indly <= P0CMDEN_indelay after IN_DELAY;
    P0CMDINSTR_indly <= P0CMDINSTR_indelay after IN_DELAY;
    P0CMDRA_indly <= P0CMDRA_indelay after IN_DELAY;
    P0RDEN_indly <= P0RDEN_indelay after IN_DELAY;
    P0RWRMASK_indly <= P0RWRMASK_indelay after IN_DELAY;
    P0WRDATA_indly <= P0WRDATA_indelay after IN_DELAY;
    P0WREN_indly <= P0WREN_indelay after IN_DELAY;
    P1ARBEN_indly <= P1ARBEN_indelay after IN_DELAY;
    P1CMDBA_indly <= P1CMDBA_indelay after IN_DELAY;
    P1CMDBL_indly <= P1CMDBL_indelay after IN_DELAY;
    P1CMDCA_indly <= P1CMDCA_indelay after IN_DELAY;
    P1CMDEN_indly <= P1CMDEN_indelay after IN_DELAY;
    P1CMDINSTR_indly <= P1CMDINSTR_indelay after IN_DELAY;
    P1CMDRA_indly <= P1CMDRA_indelay after IN_DELAY;
    P1RDEN_indly <= P1RDEN_indelay after IN_DELAY;
    P1RWRMASK_indly <= P1RWRMASK_indelay after IN_DELAY;
    P1WRDATA_indly <= P1WRDATA_indelay after IN_DELAY;
    P1WREN_indly <= P1WREN_indelay after IN_DELAY;
    P2ARBEN_indly <= P2ARBEN_indelay after IN_DELAY;
    P2CMDBA_indly <= P2CMDBA_indelay after IN_DELAY;
    P2CMDBL_indly <= P2CMDBL_indelay after IN_DELAY;
    P2CMDCA_indly <= P2CMDCA_indelay after IN_DELAY;
    P2CMDEN_indly <= P2CMDEN_indelay after IN_DELAY;
    P2CMDINSTR_indly <= P2CMDINSTR_indelay after IN_DELAY;
    P2CMDRA_indly <= P2CMDRA_indelay after IN_DELAY;
    P2EN_indly <= P2EN_indelay after IN_DELAY;
    P2WRDATA_indly <= P2WRDATA_indelay after IN_DELAY;
    P2WRMASK_indly <= P2WRMASK_indelay after IN_DELAY;
    P3ARBEN_indly <= P3ARBEN_indelay after IN_DELAY;
    P3CMDBA_indly <= P3CMDBA_indelay after IN_DELAY;
    P3CMDBL_indly <= P3CMDBL_indelay after IN_DELAY;
    P3CMDCA_indly <= P3CMDCA_indelay after IN_DELAY;
    P3CMDEN_indly <= P3CMDEN_indelay after IN_DELAY;
    P3CMDINSTR_indly <= P3CMDINSTR_indelay after IN_DELAY;
    P3CMDRA_indly <= P3CMDRA_indelay after IN_DELAY;
    P3EN_indly <= P3EN_indelay after IN_DELAY;
    P3WRDATA_indly <= P3WRDATA_indelay after IN_DELAY;
    P3WRMASK_indly <= P3WRMASK_indelay after IN_DELAY;
    P4ARBEN_indly <= P4ARBEN_indelay after IN_DELAY;
    P4CMDBA_indly <= P4CMDBA_indelay after IN_DELAY;
    P4CMDBL_indly <= P4CMDBL_indelay after IN_DELAY;
    P4CMDCA_indly <= P4CMDCA_indelay after IN_DELAY;
    P4CMDEN_indly <= P4CMDEN_indelay after IN_DELAY;
    P4CMDINSTR_indly <= P4CMDINSTR_indelay after IN_DELAY;
    P4CMDRA_indly <= P4CMDRA_indelay after IN_DELAY;
    P4EN_indly <= P4EN_indelay after IN_DELAY;
    P4WRDATA_indly <= P4WRDATA_indelay after IN_DELAY;
    P4WRMASK_indly <= P4WRMASK_indelay after IN_DELAY;
    P5ARBEN_indly <= P5ARBEN_indelay after IN_DELAY;
    P5CMDBA_indly <= P5CMDBA_indelay after IN_DELAY;
    P5CMDBL_indly <= P5CMDBL_indelay after IN_DELAY;
    P5CMDCA_indly <= P5CMDCA_indelay after IN_DELAY;
    P5CMDEN_indly <= P5CMDEN_indelay after IN_DELAY;
    P5CMDINSTR_indly <= P5CMDINSTR_indelay after IN_DELAY;
    P5CMDRA_indly <= P5CMDRA_indelay after IN_DELAY;
    P5EN_indly <= P5EN_indelay after IN_DELAY;
    P5WRDATA_indly <= P5WRDATA_indelay after IN_DELAY;
    P5WRMASK_indly <= P5WRMASK_indelay after IN_DELAY;
    PLLCE_indly <= PLLCE_indelay after IN_DELAY;
    PLLLOCK_indly <= PLLLOCK_indelay after IN_DELAY;
    RECAL_indly <= RECAL_indelay after IN_DELAY;
    SELFREFRESHENTER_indly <= SELFREFRESHENTER_indelay after IN_DELAY;
    SYSRST_indly <= SYSRST_indelay after IN_DELAY;
    UIADDR_indly <= UIADDR_indelay after IN_DELAY;
    UIADD_indly <= UIADD_indelay after IN_DELAY;
    UIBROADCAST_indly <= UIBROADCAST_indelay after IN_DELAY;
    UICMDEN_indly <= UICMDEN_indelay after IN_DELAY;
    UICMDIN_indly <= UICMDIN_indelay after IN_DELAY;
    UICMD_indly <= UICMD_indelay after IN_DELAY;
    UICS_indly <= UICS_indelay after IN_DELAY;
    UIDONECAL_indly <= UIDONECAL_indelay after IN_DELAY;
    UIDQCOUNT_indly <= UIDQCOUNT_indelay after IN_DELAY;
    UIDQLOWERDEC_indly <= UIDQLOWERDEC_indelay after IN_DELAY;
    UIDQLOWERINC_indly <= UIDQLOWERINC_indelay after IN_DELAY;
    UIDQUPPERDEC_indly <= UIDQUPPERDEC_indelay after IN_DELAY;
    UIDQUPPERINC_indly <= UIDQUPPERINC_indelay after IN_DELAY;
    UIDRPUPDATE_indly <= UIDRPUPDATE_indelay after IN_DELAY;
    UILDQSDEC_indly <= UILDQSDEC_indelay after IN_DELAY;
    UILDQSINC_indly <= UILDQSINC_indelay after IN_DELAY;
    UIREAD_indly <= UIREAD_indelay after IN_DELAY;
    UISDI_indly <= UISDI_indelay after IN_DELAY;
    UIUDQSDEC_indly <= UIUDQSDEC_indelay after IN_DELAY;
    UIUDQSINC_indly <= UIUDQSINC_indelay after IN_DELAY;
   
-- <!--Aldec correction start
	GSR_local <= GSR;
-- Aldec correction end -->

   PLLCLK_0 <= PLLCLK_dly(0); 
   PLLCLK_1 <= PLLCLK_dly(1); 
    
    MCB_INST : MCB_WRAP
      generic map (
        ARB_NUM_TIME_SLOTS   => ARB_NUM_TIME_SLOTS,
        ARB_TIME_SLOT_0      => ARB_TIME_SLOT_0_STRING,
        ARB_TIME_SLOT_1      => ARB_TIME_SLOT_1_STRING,
        ARB_TIME_SLOT_10     => ARB_TIME_SLOT_10_STRING,
        ARB_TIME_SLOT_11     => ARB_TIME_SLOT_11_STRING,
        ARB_TIME_SLOT_2      => ARB_TIME_SLOT_2_STRING,
        ARB_TIME_SLOT_3      => ARB_TIME_SLOT_3_STRING,
        ARB_TIME_SLOT_4      => ARB_TIME_SLOT_4_STRING,
        ARB_TIME_SLOT_5      => ARB_TIME_SLOT_5_STRING,
        ARB_TIME_SLOT_6      => ARB_TIME_SLOT_6_STRING,
        ARB_TIME_SLOT_7      => ARB_TIME_SLOT_7_STRING,
        ARB_TIME_SLOT_8      => ARB_TIME_SLOT_8_STRING,
        ARB_TIME_SLOT_9      => ARB_TIME_SLOT_9_STRING,
        CAL_BA               => CAL_BA_STRING,
        CAL_BYPASS           => CAL_BYPASS,
        CAL_CA               => CAL_CA_STRING,
        CAL_CALIBRATION_MODE => CAL_CALIBRATION_MODE,
        CAL_CLK_DIV          => CAL_CLK_DIV,
        CAL_DELAY            => CAL_DELAY,
        CAL_RA               => CAL_RA_STRING,
        MEM_ADDR_ORDER       => MEM_ADDR_ORDER,
        MEM_BA_SIZE          => MEM_BA_SIZE,
        MEM_BURST_LEN        => MEM_BURST_LEN,
        MEM_CAS_LATENCY      => MEM_CAS_LATENCY,
        MEM_CA_SIZE          => MEM_CA_SIZE,
        MEM_DDR1_2_ODS       => MEM_DDR1_2_ODS,
        MEM_DDR2_3_HIGH_TEMP_SR => MEM_DDR2_3_HIGH_TEMP_SR,
        MEM_DDR2_3_PA_SR     => MEM_DDR2_3_PA_SR,
        MEM_DDR2_ADD_LATENCY => MEM_DDR2_ADD_LATENCY,
        MEM_DDR2_DIFF_DQS_EN => MEM_DDR2_DIFF_DQS_EN,
        MEM_DDR2_RTT         => MEM_DDR2_RTT,
        MEM_DDR2_WRT_RECOVERY => MEM_DDR2_WRT_RECOVERY,
        MEM_DDR3_ADD_LATENCY => MEM_DDR3_ADD_LATENCY,
        MEM_DDR3_AUTO_SR     => MEM_DDR3_AUTO_SR,
        MEM_DDR3_CAS_LATENCY => MEM_DDR3_CAS_LATENCY,
        MEM_DDR3_CAS_WR_LATENCY => MEM_DDR3_CAS_WR_LATENCY,
        MEM_DDR3_DYN_WRT_ODT => MEM_DDR3_DYN_WRT_ODT,
        MEM_DDR3_ODS         => MEM_DDR3_ODS,
        MEM_DDR3_RTT         => MEM_DDR3_RTT,
        MEM_DDR3_WRT_RECOVERY => MEM_DDR3_WRT_RECOVERY,
        MEM_MDDR_ODS         => MEM_MDDR_ODS,
        MEM_MOBILE_PA_SR     => MEM_MOBILE_PA_SR,
        MEM_MOBILE_TC_SR     => MEM_MOBILE_TC_SR,
        MEM_RAS_VAL          => MEM_RAS_VAL,
        MEM_RA_SIZE          => MEM_RA_SIZE,
        MEM_RCD_VAL          => MEM_RCD_VAL,
        MEM_REFI_VAL         => MEM_REFI_VAL,
        MEM_RFC_VAL          => MEM_RFC_VAL,
        MEM_RP_VAL           => MEM_RP_VAL,
        MEM_RTP_VAL          => MEM_RTP_VAL,
        MEM_TYPE             => MEM_TYPE,
        MEM_WIDTH            => MEM_WIDTH,
        MEM_WR_VAL           => MEM_WR_VAL,
        MEM_WTR_VAL          => MEM_WTR_VAL,
        PORT_CONFIG          => PORT_CONFIG
      )
      
      port map (
        ADDR                 => ADDR_outdelay,
        BA                   => BA_outdelay,
        CAS                  => CAS_outdelay,
        CKE                  => CKE_outdelay,
        DQIOWEN0             => DQIOWEN0_outdelay,
        DQON                 => DQON_outdelay,
        DQOP                 => DQOP_outdelay,
        DQSIOWEN90N          => DQSIOWEN90N_outdelay,
        DQSIOWEN90P          => DQSIOWEN90P_outdelay,
        IOIDRPADD            => IOIDRPADD_outdelay,
        IOIDRPADDR           => IOIDRPADDR_outdelay,
        IOIDRPBROADCAST      => IOIDRPBROADCAST_outdelay,
        IOIDRPCLK            => IOIDRPCLK_outdelay,
        IOIDRPCS             => IOIDRPCS_outdelay,
        IOIDRPSDO            => IOIDRPSDO_outdelay,
        IOIDRPTRAIN          => IOIDRPTRAIN_outdelay,
        IOIDRPUPDATE         => IOIDRPUPDATE_outdelay,
        LDMN                 => LDMN_outdelay,
        LDMP                 => LDMP_outdelay,
        ODT                  => ODT_outdelay,
        P0CMDEMPTY           => P0CMDEMPTY_outdelay,
        P0CMDFULL            => P0CMDFULL_outdelay,
        P0RDCOUNT            => P0RDCOUNT_outdelay,
        P0RDDATA             => P0RDDATA_outdelay,
        P0RDEMPTY            => P0RDEMPTY_outdelay,
        P0RDERROR            => P0RDERROR_outdelay,
        P0RDFULL             => P0RDFULL_outdelay,
        P0RDOVERFLOW         => P0RDOVERFLOW_outdelay,
        P0WRCOUNT            => P0WRCOUNT_outdelay,
        P0WREMPTY            => P0WREMPTY_outdelay,
        P0WRERROR            => P0WRERROR_outdelay,
        P0WRFULL             => P0WRFULL_outdelay,
        P0WRUNDERRUN         => P0WRUNDERRUN_outdelay,
        P1CMDEMPTY           => P1CMDEMPTY_outdelay,
        P1CMDFULL            => P1CMDFULL_outdelay,
        P1RDCOUNT            => P1RDCOUNT_outdelay,
        P1RDDATA             => P1RDDATA_outdelay,
        P1RDEMPTY            => P1RDEMPTY_outdelay,
        P1RDERROR            => P1RDERROR_outdelay,
        P1RDFULL             => P1RDFULL_outdelay,
        P1RDOVERFLOW         => P1RDOVERFLOW_outdelay,
        P1WRCOUNT            => P1WRCOUNT_outdelay,
        P1WREMPTY            => P1WREMPTY_outdelay,
        P1WRERROR            => P1WRERROR_outdelay,
        P1WRFULL             => P1WRFULL_outdelay,
        P1WRUNDERRUN         => P1WRUNDERRUN_outdelay,
        P2CMDEMPTY           => P2CMDEMPTY_outdelay,
        P2CMDFULL            => P2CMDFULL_outdelay,
        P2COUNT              => P2COUNT_outdelay,
        P2EMPTY              => P2EMPTY_outdelay,
        P2ERROR              => P2ERROR_outdelay,
        P2FULL               => P2FULL_outdelay,
        P2RDDATA             => P2RDDATA_outdelay,
        P2RDOVERFLOW         => P2RDOVERFLOW_outdelay,
        P2WRUNDERRUN         => P2WRUNDERRUN_outdelay,
        P3CMDEMPTY           => P3CMDEMPTY_outdelay,
        P3CMDFULL            => P3CMDFULL_outdelay,
        P3COUNT              => P3COUNT_outdelay,
        P3EMPTY              => P3EMPTY_outdelay,
        P3ERROR              => P3ERROR_outdelay,
        P3FULL               => P3FULL_outdelay,
        P3RDDATA             => P3RDDATA_outdelay,
        P3RDOVERFLOW         => P3RDOVERFLOW_outdelay,
        P3WRUNDERRUN         => P3WRUNDERRUN_outdelay,
        P4CMDEMPTY           => P4CMDEMPTY_outdelay,
        P4CMDFULL            => P4CMDFULL_outdelay,
        P4COUNT              => P4COUNT_outdelay,
        P4EMPTY              => P4EMPTY_outdelay,
        P4ERROR              => P4ERROR_outdelay,
        P4FULL               => P4FULL_outdelay,
        P4RDDATA             => P4RDDATA_outdelay,
        P4RDOVERFLOW         => P4RDOVERFLOW_outdelay,
        P4WRUNDERRUN         => P4WRUNDERRUN_outdelay,
        P5CMDEMPTY           => P5CMDEMPTY_outdelay,
        P5CMDFULL            => P5CMDFULL_outdelay,
        P5COUNT              => P5COUNT_outdelay,
        P5EMPTY              => P5EMPTY_outdelay,
        P5ERROR              => P5ERROR_outdelay,
        P5FULL               => P5FULL_outdelay,
        P5RDDATA             => P5RDDATA_outdelay,
        P5RDOVERFLOW         => P5RDOVERFLOW_outdelay,
        P5WRUNDERRUN         => P5WRUNDERRUN_outdelay,
        RAS                  => RAS_outdelay,
        RST                  => RST_outdelay,
        SELFREFRESHMODE      => SELFREFRESHMODE_outdelay,
        STATUS               => STATUS_outdelay,
        UDMN                 => UDMN_outdelay,
        UDMP                 => UDMP_outdelay,
        UOCALSTART           => UOCALSTART_outdelay,
        UOCMDREADYIN         => UOCMDREADYIN_outdelay,
        UODATA               => UODATA_outdelay,
        UODATAVALID          => UODATAVALID_outdelay,
        UODONECAL            => UODONECAL_outdelay,
        UOREFRSHFLAG         => UOREFRSHFLAG_outdelay,
        UOSDO                => UOSDO_outdelay,
        WE                   => WE_outdelay,
        DQI                  => DQI_indly,
        DQSIOIN              => DQSIOIN_indly,
        DQSIOIP              => DQSIOIP_indly,
        IOIDRPSDI            => IOIDRPSDI_indly,
        P0ARBEN              => P0ARBEN_indly,
        P0CMDBA              => P0CMDBA_indly,
        P0CMDBL              => P0CMDBL_indly,
        P0CMDCA              => P0CMDCA_indly,
        P0CMDCLK             => P0CMDCLK_indly,
        P0CMDEN              => P0CMDEN_indly,
        P0CMDINSTR           => P0CMDINSTR_indly,
        P0CMDRA              => P0CMDRA_indly,
        P0RDCLK              => P0RDCLK_indly,
        P0RDEN               => P0RDEN_indly,
        P0RWRMASK            => P0RWRMASK_indly,
        P0WRCLK              => P0WRCLK_indly,
        P0WRDATA             => P0WRDATA_indly,
        P0WREN               => P0WREN_indly,
        P1ARBEN              => P1ARBEN_indly,
        P1CMDBA              => P1CMDBA_indly,
        P1CMDBL              => P1CMDBL_indly,
        P1CMDCA              => P1CMDCA_indly,
        P1CMDCLK             => P1CMDCLK_indly,
        P1CMDEN              => P1CMDEN_indly,
        P1CMDINSTR           => P1CMDINSTR_indly,
        P1CMDRA              => P1CMDRA_indly,
        P1RDCLK              => P1RDCLK_indly,
        P1RDEN               => P1RDEN_indly,
        P1RWRMASK            => P1RWRMASK_indly,
        P1WRCLK              => P1WRCLK_indly,
        P1WRDATA             => P1WRDATA_indly,
        P1WREN               => P1WREN_indly,
        P2ARBEN              => P2ARBEN_indly,
        P2CLK                => P2CLK_indly,
        P2CMDBA              => P2CMDBA_indly,
        P2CMDBL              => P2CMDBL_indly,
        P2CMDCA              => P2CMDCA_indly,
        P2CMDCLK             => P2CMDCLK_indly,
        P2CMDEN              => P2CMDEN_indly,
        P2CMDINSTR           => P2CMDINSTR_indly,
        P2CMDRA              => P2CMDRA_indly,
        P2EN                 => P2EN_indly,
        P2WRDATA             => P2WRDATA_indly,
        P2WRMASK             => P2WRMASK_indly,
        P3ARBEN              => P3ARBEN_indly,
        P3CLK                => P3CLK_indly,
        P3CMDBA              => P3CMDBA_indly,
        P3CMDBL              => P3CMDBL_indly,
        P3CMDCA              => P3CMDCA_indly,
        P3CMDCLK             => P3CMDCLK_indly,
        P3CMDEN              => P3CMDEN_indly,
        P3CMDINSTR           => P3CMDINSTR_indly,
        P3CMDRA              => P3CMDRA_indly,
        P3EN                 => P3EN_indly,
        P3WRDATA             => P3WRDATA_indly,
        P3WRMASK             => P3WRMASK_indly,
        P4ARBEN              => P4ARBEN_indly,
        P4CLK                => P4CLK_indly,
        P4CMDBA              => P4CMDBA_indly,
        P4CMDBL              => P4CMDBL_indly,
        P4CMDCA              => P4CMDCA_indly,
        P4CMDCLK             => P4CMDCLK_indly,
        P4CMDEN              => P4CMDEN_indly,
        P4CMDINSTR           => P4CMDINSTR_indly,
        P4CMDRA              => P4CMDRA_indly,
        P4EN                 => P4EN_indly,
        P4WRDATA             => P4WRDATA_indly,
        P4WRMASK             => P4WRMASK_indly,
        P5ARBEN              => P5ARBEN_indly,
        P5CLK                => P5CLK_indly,
        P5CMDBA              => P5CMDBA_indly,
        P5CMDBL              => P5CMDBL_indly,
        P5CMDCA              => P5CMDCA_indly,
        P5CMDCLK             => P5CMDCLK_indly,
        P5CMDEN              => P5CMDEN_indly,
        P5CMDINSTR           => P5CMDINSTR_indly,
        P5CMDRA              => P5CMDRA_indly,
        P5EN                 => P5EN_indly,
        P5WRDATA             => P5WRDATA_indly,
        P5WRMASK             => P5WRMASK_indly,
        PLLCE                => PLLCE_indly,
        PLLCLK               => PLLCLK_indly,
        PLLLOCK              => PLLLOCK_indly,
        RECAL                => RECAL_indly,
        SELFREFRESHENTER     => SELFREFRESHENTER_indly,
        SYSRST               => SYSRST_indly,
        UDQSIOIN             => UDQSIOIN_indly,
        UDQSIOIP             => UDQSIOIP_indly,
        UIADD                => UIADD_indly,
        UIADDR               => UIADDR_indly,
        UIBROADCAST          => UIBROADCAST_indly,
        UICLK                => UICLK_indly,
        UICMD                => UICMD_indly,
        UICMDEN              => UICMDEN_indly,
        UICMDIN              => UICMDIN_indly,
        UICS                 => UICS_indly,
        UIDONECAL            => UIDONECAL_indly,
        UIDQCOUNT            => UIDQCOUNT_indly,
        UIDQLOWERDEC         => UIDQLOWERDEC_indly,
        UIDQLOWERINC         => UIDQLOWERINC_indly,
        UIDQUPPERDEC         => UIDQUPPERDEC_indly,
        UIDQUPPERINC         => UIDQUPPERINC_indly,
        UIDRPUPDATE          => UIDRPUPDATE_indly,
        UILDQSDEC            => UILDQSDEC_indly,
        UILDQSINC            => UILDQSINC_indly,
        UIREAD               => UIREAD_indly,
        UISDI                => UISDI_indly,
        UIUDQSDEC            => UIUDQSDEC_indly,
        UIUDQSINC            => UIUDQSINC_indly,        
-- <!--Aldec correction start        
        GSR => GSR_local
-- Aldec correction end -->
      );
    
    INIPROC : process
    begin
      -- case CAL_BYPASS is
      if((CAL_BYPASS = "YES") or (CAL_BYPASS = "yes")) then
        CAL_BYPASS_BINARY <= '1';
      elsif((CAL_BYPASS = "NO") or (CAL_BYPASS= "no")) then
        CAL_BYPASS_BINARY <= '0';
      else
        assert FALSE report "Error : CAL_BYPASS = is not YES, NO." severity error;
      end if;
    -- end case;
    -- case CAL_CALIBRATION_MODE is
      if((CAL_CALIBRATION_MODE = "CALIBRATION") or (CAL_CALIBRATION_MODE = "calibration")) then
        CAL_CALIBRATION_MODE_BINARY <= '0';
      elsif((CAL_CALIBRATION_MODE = "NOCALIBRATION") or (CAL_CALIBRATION_MODE= "nocalibration")) then
        CAL_CALIBRATION_MODE_BINARY <= '1';
      else
        assert FALSE report "Error : CAL_CALIBRATION_MODE = is not CALIBRATION, NOCALIBRATION." severity error;
      end if;
    -- end case;
    -- case CAL_DELAY is
      if((CAL_DELAY = "QUARTER") or (CAL_DELAY = "quarter")) then
        CAL_DELAY_BINARY <= "00";
      elsif((CAL_DELAY = "FULL") or (CAL_DELAY= "full")) then
        CAL_DELAY_BINARY <= "11";
      elsif((CAL_DELAY = "HALF") or (CAL_DELAY= "half")) then
        CAL_DELAY_BINARY <= "01";
      elsif((CAL_DELAY = "THREEQUARTER") or (CAL_DELAY= "threequarter")) then
        CAL_DELAY_BINARY <= "10";
      else
        assert FALSE report "Error : CAL_DELAY = is not QUARTER, FULL, HALF, THREEQUARTER." severity error;
      end if;
    -- end case;
     -- case MEM_TYPE is
      if((MEM_TYPE = "DDR3") or (MEM_TYPE = "ddr3")) then
        MEM_TYPE_BINARY <= "000";
      elsif((MEM_TYPE = "DDR") or (MEM_TYPE= "ddr")) then
        MEM_TYPE_BINARY <= "010";
      elsif((MEM_TYPE = "DDR2") or (MEM_TYPE= "ddr2")) then
        MEM_TYPE_BINARY <= "001";
      elsif((MEM_TYPE = "MDDR") or (MEM_TYPE= "mddr")) then
        MEM_TYPE_BINARY <= "011";
      else
        assert FALSE report "Error : MEM_TYPE = is not DDR3, DDR, DDR2, MDDR." severity error;
      end if;
    -- end case;
    -- case MEM_BURST_LEN is
     if (MEM_BURST_LEN = 4)  then
      if (MEM_TYPE = "DDR3") then
        assert FALSE report "Error : MEM_BURST_LEN of 4 is not allowed for MEM_TYPE DDR3." severity error;
      else
        MEM_BURST_LEN_BINARY <= "010";
      end if;
     elsif (MEM_BURST_LEN = 8) then
      MEM_BURST_LEN_BINARY <= "011";
     else
      assert FALSE report "Error : MEM_BURST_LEN is not 4 or 8." severity error;
     end if;
    -- end case
    -- case MEM_ADDR_ORDER is
      if((MEM_ADDR_ORDER = "BANK_ROW_COLUMN") or (MEM_ADDR_ORDER = "bank_row_column")) then
        MEM_ADDR_ORDER_BINARY <= '0';
      elsif((MEM_ADDR_ORDER = "ROW_BANK_COLUMN") or (MEM_ADDR_ORDER= "row_bank_column")) then
        MEM_ADDR_ORDER_BINARY <= '1';
      else
        assert FALSE report "Error : MEM_ADDR_ORDER = is not BANK_ROW_COLUMN, ROW_BANK_COLUMN." severity error;
      end if;
    -- end case;
    -- case MEM_DDR1_2_ODS is
    if ((MEM_TYPE = "DDR2") or (MEM_TYPE = "DDR")) then
      if((MEM_DDR1_2_ODS = "FULL") or (MEM_DDR1_2_ODS = "full")) then
        MEM_DDR1_2_ODS_BINARY <= '0';
      elsif((MEM_DDR1_2_ODS = "REDUCED") or (MEM_DDR1_2_ODS= "reduced")) then
        MEM_DDR1_2_ODS_BINARY <= '1';
      else
        assert FALSE report "Error : MEM_DDR1_2_ODS = is not FULL, REDUCED." severity error;
      end if;
    end if;
    -- end case;
    -- case MEM_DDR2_3_HIGH_TEMP_SR is
    if ((MEM_TYPE = "DDR2") or (MEM_TYPE = "DDR3")) then
      if((MEM_DDR2_3_HIGH_TEMP_SR = "NORMAL") or (MEM_DDR2_3_HIGH_TEMP_SR = "normal")) then
        MEM_DDR2_3_HIGH_TEMP_SR_BINARY <= '0';
      elsif((MEM_DDR2_3_HIGH_TEMP_SR = "EXTENDED") or (MEM_DDR2_3_HIGH_TEMP_SR= "extended")) then
        MEM_DDR2_3_HIGH_TEMP_SR_BINARY <= '1';
      else
        assert FALSE report "Error : MEM_DDR2_3_HIGH_TEMP_SR = is not NORMAL, EXTENDED." severity error;
      end if;
    -- end case;
    -- case MEM_DDR2_3_PA_SR is
      if((MEM_DDR2_3_PA_SR = "FULL") or (MEM_DDR2_3_PA_SR = "full")) then
        MEM_DDR2_3_PA_SR_BINARY <= "000";
      elsif((MEM_DDR2_3_PA_SR = "EIGHTH1") or (MEM_DDR2_3_PA_SR= "eighth1")) then
        MEM_DDR2_3_PA_SR_BINARY <= "011";
      elsif((MEM_DDR2_3_PA_SR = "EIGHTH2") or (MEM_DDR2_3_PA_SR= "eighth2")) then
        MEM_DDR2_3_PA_SR_BINARY <= "111";
      elsif((MEM_DDR2_3_PA_SR = "HALF1") or (MEM_DDR2_3_PA_SR= "half1")) then
        MEM_DDR2_3_PA_SR_BINARY <= "001";
      elsif((MEM_DDR2_3_PA_SR = "HALF2") or (MEM_DDR2_3_PA_SR= "half2")) then
        MEM_DDR2_3_PA_SR_BINARY <= "101";
      elsif((MEM_DDR2_3_PA_SR = "QUARTER1") or (MEM_DDR2_3_PA_SR= "quarter1")) then
        MEM_DDR2_3_PA_SR_BINARY <= "010";
      elsif((MEM_DDR2_3_PA_SR = "QUARTER2") or (MEM_DDR2_3_PA_SR= "quarter2")) then
        MEM_DDR2_3_PA_SR_BINARY <= "110";
      elsif((MEM_DDR2_3_PA_SR = "THREEQUARTER") or (MEM_DDR2_3_PA_SR= "threequarter")) then
        MEM_DDR2_3_PA_SR_BINARY <= "100";
      else
        assert FALSE report "Error : MEM_DDR2_3_PA_SR = is not FULL, EIGHTH1, EIGHTH2, HALF1, HALF2, QUARTER1, QUARTER2, THREEQUARTER." severity error;
      end if;
    end if;
    -- end case;
    -- case MEM_DDR2_DIFF_DQS_EN is
    if (MEM_TYPE = "DDR2") then
      if((MEM_DDR2_DIFF_DQS_EN = "YES") or (MEM_DDR2_DIFF_DQS_EN = "yes")) then
        MEM_DDR2_DIFF_DQS_EN_BINARY <= '0';
      elsif((MEM_DDR2_DIFF_DQS_EN = "NO") or (MEM_DDR2_DIFF_DQS_EN= "no")) then
        MEM_DDR2_DIFF_DQS_EN_BINARY <= '1';
      else
        assert FALSE report "Error : MEM_DDR2_DIFF_DQS_EN = is not YES, NO." severity error;
      end if;
    -- end case;
    -- case MEM_DDR2_RTT is
      if((MEM_DDR2_RTT = "50OHMS") or (MEM_DDR2_RTT = "50ohms")) then
        MEM_DDR2_RTT_BINARY <= "11";
      elsif((MEM_DDR2_RTT = "75OHMS") or (MEM_DDR2_RTT= "75ohms")) then
        MEM_DDR2_RTT_BINARY <= "01";
      elsif((MEM_DDR2_RTT = "150OHMS") or (MEM_DDR2_RTT= "150ohms")) then
        MEM_DDR2_RTT_BINARY <= "10";
      elsif((MEM_DDR2_RTT = "OFF") or (MEM_DDR2_RTT= "off")) then
        MEM_DDR2_RTT_BINARY <= "00";
      else
        assert FALSE report "Error : MEM_DDR2_RTT = is not 50OHMS, 75OHMS, 150OHMS, OFF." severity error;
      end if;
      if ((MEM_DDR2_ADD_LATENCY >= 0) and (MEM_DDR2_ADD_LATENCY <= 5)) then
        MEM_DDR2_ADD_LATENCY_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_DDR2_ADD_LATENCY, 3);
      else
       assert FALSE report "Error : MEM_DDR2_ADD_LATENCY is not in range 0 .. 5." severity error;
      end if;
      if ((MEM_DDR2_WRT_RECOVERY >= 2) and (MEM_DDR2_WRT_RECOVERY <= 6)) then
        MEM_DDR2_WRT_RECOVERY_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_DDR2_WRT_RECOVERY, 3);
      else
       assert FALSE report "Error : MEM_DDR2_WRT_RECOVERY is not in range 2 .. 6." severity error;
      end if;

    end if;
    -- end case;
    -- case MEM_DDR3_ADD_LATENCY is
    if (MEM_TYPE = "DDR3") then
      if((MEM_DDR3_ADD_LATENCY = "OFF") or (MEM_DDR3_ADD_LATENCY = "off")) then
        MEM_DDR3_ADD_LATENCY_BINARY <= "00";
      elsif((MEM_DDR3_ADD_LATENCY = "CL1") or (MEM_DDR3_ADD_LATENCY= "cl1")) then
        MEM_DDR3_ADD_LATENCY_BINARY <= "01";
      elsif((MEM_DDR3_ADD_LATENCY = "CL2") or (MEM_DDR3_ADD_LATENCY= "cl2")) then
        MEM_DDR3_ADD_LATENCY_BINARY <= "10";
      else
        assert FALSE report "Error : MEM_DDR3_ADD_LATENCY = is not OFF, CL1, CL2." severity error;
      end if;
    -- end case;
    -- case MEM_DDR3_AUTO_SR is
      if((MEM_DDR3_AUTO_SR = "ENABLED") or (MEM_DDR3_AUTO_SR = "enabled")) then
        MEM_DDR3_AUTO_SR_BINARY <= '1';
      elsif((MEM_DDR3_AUTO_SR = "MANUAL") or (MEM_DDR3_AUTO_SR= "manual")) then
        MEM_DDR3_AUTO_SR_BINARY <= '0';
      else
        assert FALSE report "Error : MEM_DDR3_AUTO_SR = is not ENABLED, MANUAL." severity error;
      end if;
    -- end case;
    -- case MEM_DDR3_DYN_WRT_ODT is
      if((MEM_DDR3_DYN_WRT_ODT = "OFF") or (MEM_DDR3_DYN_WRT_ODT = "off")) then
        MEM_DDR3_DYN_WRT_ODT_BINARY <= "00";
      elsif((MEM_DDR3_DYN_WRT_ODT = "DIV2") or (MEM_DDR3_DYN_WRT_ODT= "div2")) then
        MEM_DDR3_DYN_WRT_ODT_BINARY <= "01";
      elsif((MEM_DDR3_DYN_WRT_ODT = "DIV4") or (MEM_DDR3_DYN_WRT_ODT= "div4")) then
        MEM_DDR3_DYN_WRT_ODT_BINARY <= "10";
      else
        assert FALSE report "Error : MEM_DDR3_DYN_WRT_ODT = is not OFF, DIV2, DIV4." severity error;
      end if;
    -- end case;
    -- case MEM_DDR3_ODS is
      if((MEM_DDR3_ODS = "DIV7") or (MEM_DDR3_ODS = "div7")) then
        MEM_DDR3_ODS_BINARY <= "01";
      elsif((MEM_DDR3_ODS = "DIV6") or (MEM_DDR3_ODS= "div6")) then
        MEM_DDR3_ODS_BINARY <= "00";
      else
        assert FALSE report "Error : MEM_DDR3_ODS = is not DIV7, DIV6." severity error;
      end if;
    -- end case;
    -- case MEM_DDR3_RTT is
      if((MEM_DDR3_RTT = "DIV2") or (MEM_DDR3_RTT = "div2")) then
        MEM_DDR3_RTT_BINARY <= "010";
      elsif((MEM_DDR3_RTT = "DIV4") or (MEM_DDR3_RTT= "div4")) then
        MEM_DDR3_RTT_BINARY <= "001";
      elsif((MEM_DDR3_RTT = "DIV6") or (MEM_DDR3_RTT= "div6")) then
        MEM_DDR3_RTT_BINARY <= "011";
      elsif((MEM_DDR3_RTT = "DIV8") or (MEM_DDR3_RTT= "div8")) then
        MEM_DDR3_RTT_BINARY <= "100";
      elsif((MEM_DDR3_RTT = "DIV12") or (MEM_DDR3_RTT= "div12")) then
        MEM_DDR3_RTT_BINARY <= "101";
      elsif((MEM_DDR3_RTT = "OFF") or (MEM_DDR3_RTT= "off")) then
        MEM_DDR3_RTT_BINARY <= "000";
      else
        assert FALSE report "Error : MEM_DDR3_RTT = is not DIV2, DIV4, DIV6, DIV8, DIV12, OFF." severity error;
      end if;
      if ((MEM_DDR3_CAS_LATENCY >= 5) and (MEM_DDR3_CAS_LATENCY <= 10)) then
      MEM_DDR3_CAS_LATENCY_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_DDR3_CAS_LATENCY, 4);
      else
        assert FALSE report "Error : MEM_DDR3_CAS_LATENCY is not in range 5 .. 10." severity error;
      end if;
      if ((MEM_DDR3_CAS_WR_LATENCY >= 5) and (MEM_DDR3_CAS_WR_LATENCY <= 8)) then
       MEM_DDR3_CAS_WR_LATENCY_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_DDR3_CAS_WR_LATENCY, 3);
      else
        assert FALSE report "Error : MEM_DDR3_CAS_WR_LATENCY is not in range 5 .. 8." severity error;
      end if;
      if ((MEM_DDR3_WRT_RECOVERY = 5) or (MEM_DDR3_WRT_RECOVERY = 6) or (MEM_DDR3_WRT_RECOVERY = 7) or (MEM_DDR3_WRT_RECOVERY = 8) or (MEM_DDR3_WRT_RECOVERY = 10) or (MEM_DDR3_WRT_RECOVERY = 12)) then
        MEM_DDR3_WRT_RECOVERY_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_DDR3_WRT_RECOVERY, 3);
      else
       assert FALSE report "Error : MEM_DDR3_WRT_RECOVERY is not 5, 6, 7, 8, 10 or 12." severity error;
      end if;
    end if;
    -- end case;
    -- case MEM_MDDR_ODS is
    if (MEM_TYPE = "MDDR") then
      if((MEM_MDDR_ODS = "FULL") or (MEM_MDDR_ODS = "full")) then
        MEM_MDDR_ODS_BINARY <= "000";
      elsif((MEM_MDDR_ODS = "HALF") or (MEM_MDDR_ODS= "half")) then
        MEM_MDDR_ODS_BINARY <= "001";
      elsif((MEM_MDDR_ODS = "QUARTER") or (MEM_MDDR_ODS= "quarter")) then
        MEM_MDDR_ODS_BINARY <= "010";
      elsif((MEM_MDDR_ODS = "THREEQUARTERS") or (MEM_MDDR_ODS= "threequarters")) then
        MEM_MDDR_ODS_BINARY <= "100";
      else
        assert FALSE report "Error : MEM_MDDR_ODS = is not FULL, HALF, QUARTER, THREEQUARTERS." severity error;
      end if;
    -- end case;
    -- case MEM_MOBILE_PA_SR is
      if((MEM_MOBILE_PA_SR = "FULL") or (MEM_MOBILE_PA_SR = "full")) then
        MEM_MOBILE_PA_SR_BINARY <= "000";
      elsif((MEM_MOBILE_PA_SR = "HALF") or (MEM_MOBILE_PA_SR= "half")) then
        MEM_MOBILE_PA_SR_BINARY <= "001";
      else
        assert FALSE report "Error : MEM_MOBILE_PA_SR = is not FULL, HALF." severity error;
      end if;
       if ((MEM_MOBILE_TC_SR >= 0) and (MEM_MOBILE_TC_SR <= 3)) then
        MEM_MOBILE_TC_SR_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_MOBILE_TC_SR, 2);
       else
        assert FALSE report "Error : MEM_MOBILE_TC_SR is not in range 0 .. 3." severity error;
      end if;
     end if;
    -- end case;
    case ARB_NUM_TIME_SLOTS is
      when  12   =>  ARB_NUM_TIME_SLOTS_BINARY <= '1';
      when  10   =>  ARB_NUM_TIME_SLOTS_BINARY <= '0';
      when others  =>  assert FALSE report "Error : ARB_NUM_TIME_SLOTS is 12 or 10." severity error;
    end case;
    case MEM_BA_SIZE is
      when  3   =>  MEM_BA_SIZE_BINARY <= '1';
      when  2   =>  MEM_BA_SIZE_BINARY <= '0';
      when others  =>  assert FALSE report "Error : MEM_BA_SIZE is not in range 2 .. 3." severity error;
    end case;
    if ((CAL_CLK_DIV = 1) or (CAL_CLK_DIV = 2) or (CAL_CLK_DIV = 4) or (CAL_CLK_DIV = 8)) then
      CAL_CLK_DIV_BINARY <= CONV_STD_LOGIC_VECTOR(CAL_CLK_DIV, 3);
    else
      assert FALSE report "Error : CAL_CLK_DIV is not  1, 2, 4 or 8." severity error;
    end if;
    if ((MEM_CAS_LATENCY >= 1) and (MEM_CAS_LATENCY <= 6)) then
      MEM_CAS_LATENCY_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_CAS_LATENCY, 3);
    else
      assert FALSE report "Error : MEM_CAS_LATENCY is not in range 1 .. 6." severity error;
    end if;
    if ((MEM_CA_SIZE >= 9) and (MEM_CA_SIZE <= 12)) then
      MEM_CA_SIZE_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_CA_SIZE, 2);
    else
      assert FALSE report "Error : MEM_CA_SIZE is not in range 9 .. 12." severity error;
    end if;
    if ((MEM_RAS_VAL >= 0) and (MEM_RAS_VAL <= 31)) then
      MEM_RAS_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_RAS_VAL, 5);
    else
      assert FALSE report "Error : MEM_RAS_VAL is not in range 0 .. 31." severity error;
    end if;
    if ((MEM_RA_SIZE >= 12) and (MEM_RA_SIZE <= 15)) then
      MEM_RA_SIZE_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_RA_SIZE, 2);
    else
      assert FALSE report "Error : MEM_RA_SIZE is not in range 12 .. 15." severity error;
    end if;
    if ((MEM_RCD_VAL >= 0) and (MEM_RCD_VAL <= 7)) then
      MEM_RCD_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_RCD_VAL, 3);
    else
      assert FALSE report "Error : MEM_RCD_VAL is not in range 0 .. 7." severity error;
    end if;
    if ((MEM_REFI_VAL >= 0) and (MEM_REFI_VAL <= 4095)) then
      MEM_REFI_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_REFI_VAL, 12);
    else
      assert FALSE report "Error : MEM_REFI_VAL is not in range 0 .. 4095." severity error;
    end if;
    if ((MEM_RFC_VAL >= 0) and (MEM_RFC_VAL <= 255)) then
      MEM_RFC_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_RFC_VAL, 8);
    else
      assert FALSE report "Error : MEM_RFC_VAL is not in range 0 .. 255." severity error;
    end if;
    if ((MEM_RP_VAL >= 0) and (MEM_RP_VAL <= 15)) then
      MEM_RP_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_RP_VAL, 4);
    else
      assert FALSE report "Error : MEM_RP_VAL is not in range 0 .. 15." severity error;
    end if;
    if ((MEM_RTP_VAL >= 0) and (MEM_RTP_VAL <= 7)) then
      MEM_RTP_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_RTP_VAL, 3);
    else
      assert FALSE report "Error : MEM_RTP_VAL is not in range 0 .. 7." severity error;
    end if;
    if ((MEM_WIDTH = 4) or (MEM_WIDTH = 8) or (MEM_WIDTH = 16)) then
      MEM_WIDTH_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_WIDTH, 2);
    else
      assert FALSE report "Error : MEM_WIDTH is not 4, 8 or 16." severity error;
    end if;
    if ((MEM_WR_VAL >= 0) and (MEM_WR_VAL <= 7)) then
      MEM_WR_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_WR_VAL, 3);
    else
      assert FALSE report "Error : MEM_WR_VAL is not in range 0 .. 7." severity error;
    end if;
    if ((MEM_WTR_VAL >= 0) and (MEM_WTR_VAL <= 7)) then
      MEM_WTR_VAL_BINARY <= CONV_STD_LOGIC_VECTOR(MEM_WTR_VAL, 3);
    else
      assert FALSE report "Error : MEM_WTR_VAL is not in range 0 .. 7." severity error;
    end if;
     -- case PORT_CONFIG is
      if((PORT_CONFIG = "B32_B32_B32_B32") or (PORT_CONFIG = "b32_b32_b32_b32")) then
        PORT_CONFIG_BINARY <= "001";
      elsif((PORT_CONFIG = "B32_B32_R32_R32_R32_R32") or (PORT_CONFIG= "b32_b32_r32_r32_r32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_R32_R32_W32") or (PORT_CONFIG= "b32_b32_r32_r32_r32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_R32_W32_R32") or (PORT_CONFIG= "b32_b32_r32_r32_w32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_R32_W32_W32") or (PORT_CONFIG= "b32_b32_r32_r32_w32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_W32_R32_R32") or (PORT_CONFIG= "b32_b32_r32_w32_r32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_W32_R32_W32") or (PORT_CONFIG= "b32_b32_r32_w32_r32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_W32_W32_R32") or (PORT_CONFIG= "b32_b32_r32_w32_w32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_R32_W32_W32_W32") or (PORT_CONFIG= "b32_b32_r32_w32_w32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_R32_R32_R32") or (PORT_CONFIG= "b32_b32_w32_r32_r32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_R32_R32_W32") or (PORT_CONFIG= "b32_b32_w32_r32_r32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_R32_W32_R32") or (PORT_CONFIG= "b32_b32_w32_r32_w32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_R32_W32_W32") or (PORT_CONFIG= "b32_b32_w32_r32_w32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_W32_R32_R32") or (PORT_CONFIG= "b32_b32_w32_w32_r32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_W32_R32_W32") or (PORT_CONFIG= "b32_b32_w32_w32_r32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_W32_W32_R32") or (PORT_CONFIG= "b32_b32_w32_w32_w32_r32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B32_B32_W32_W32_W32_W32") or (PORT_CONFIG= "b32_b32_w32_w32_w32_w32")) then
        PORT_CONFIG_BINARY <= "000";
      elsif((PORT_CONFIG = "B64_B32_B32") or (PORT_CONFIG= "b64_b32_b32")) then
        PORT_CONFIG_BINARY <= "010";
      elsif((PORT_CONFIG = "B64_B64") or (PORT_CONFIG= "b64_b64")) then
        PORT_CONFIG_BINARY <= "011";
      elsif((PORT_CONFIG = "B128") or (PORT_CONFIG= "b128")) then
        PORT_CONFIG_BINARY <= "100";
      else
        assert FALSE report "Error : PORT_CONFIG = is not B32_B32_B32_B32, B32_B32_R32_R32_R32_R32, B32_B32_R32_R32_R32_W32, B32_B32_R32_R32_W32_R32, B32_B32_R32_R32_W32_W32, B32_B32_R32_W32_R32_R32, B32_B32_R32_W32_R32_W32, B32_B32_R32_W32_W32_R32, B32_B32_R32_W32_W32_W32, B32_B32_W32_R32_R32_R32, B32_B32_W32_R32_R32_W32, B32_B32_W32_R32_W32_R32, B32_B32_W32_R32_W32_W32, B32_B32_W32_W32_R32_R32, B32_B32_W32_W32_R32_W32, B32_B32_W32_W32_W32_R32, B32_B32_W32_W32_W32_W32, B64_B32_B32, B64_B64, B128." severity error;
      end if;
    -- end case;
      wait;
    end process INIPROC;
    
    TIMING : process
      variable Tmkr_IOIDRPSDI_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P0ARBEN_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_P0ARBEN_PLLCLK_0_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P0ARBEN_PLLCLK_1_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P0CMDBA_P0CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P0CMDBL_P0CMDCLK_posedge : VitalTimingDataArrayType(5 downto 0);
      variable Tmkr_P0CMDCA_P0CMDCLK_posedge : VitalTimingDataArrayType(11 downto 0);
      variable Tmkr_P0CMDEN_P0CMDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P0CMDINSTR_P0CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P0CMDRA_P0CMDCLK_posedge : VitalTimingDataArrayType(14 downto 0);
      variable Tmkr_P0RDEN_P0RDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P0RWRMASK_P0WRCLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_P0WRDATA_P0WRCLK_posedge : VitalTimingDataArrayType(31 downto 0);
      variable Tmkr_P0WREN_P0WRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P1ARBEN_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_P1CMDBA_P1CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P1CMDBL_P1CMDCLK_posedge : VitalTimingDataArrayType(5 downto 0);
      variable Tmkr_P1CMDCA_P1CMDCLK_posedge : VitalTimingDataArrayType(11 downto 0);
      variable Tmkr_P1CMDEN_P1CMDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P1CMDINSTR_P1CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P1CMDRA_P1CMDCLK_posedge : VitalTimingDataArrayType(14 downto 0);
      variable Tmkr_P1RDEN_P1RDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P1RWRMASK_P1WRCLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_P1WRDATA_P1WRCLK_posedge : VitalTimingDataArrayType(31 downto 0);
      variable Tmkr_P1WREN_P1WRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P2ARBEN_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_P2CMDBA_P2CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P2CMDBL_P2CMDCLK_posedge : VitalTimingDataArrayType(5 downto 0);
      variable Tmkr_P2CMDCA_P2CMDCLK_posedge : VitalTimingDataArrayType(11 downto 0);
      variable Tmkr_P2CMDEN_P2CMDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P2CMDINSTR_P2CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P2CMDRA_P2CMDCLK_posedge : VitalTimingDataArrayType(14 downto 0);
      variable Tmkr_P2EN_P2CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P2WRDATA_P2CLK_posedge : VitalTimingDataArrayType(31 downto 0);
      variable Tmkr_P2WRMASK_P2CLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_P3ARBEN_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_P3CMDBA_P3CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P3CMDBL_P3CMDCLK_posedge : VitalTimingDataArrayType(5 downto 0);
      variable Tmkr_P3CMDCA_P3CMDCLK_posedge : VitalTimingDataArrayType(11 downto 0);
      variable Tmkr_P3CMDEN_P3CMDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P3CMDINSTR_P3CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P3CMDRA_P3CMDCLK_posedge : VitalTimingDataArrayType(14 downto 0);
      variable Tmkr_P3EN_P3CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P3WRDATA_P3CLK_posedge : VitalTimingDataArrayType(31 downto 0);
      variable Tmkr_P3WRMASK_P3CLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_P4ARBEN_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_P4CMDBA_P4CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P4CMDBL_P4CMDCLK_posedge : VitalTimingDataArrayType(5 downto 0);
      variable Tmkr_P4CMDCA_P4CMDCLK_posedge : VitalTimingDataArrayType(11 downto 0);
      variable Tmkr_P4CMDEN_P4CMDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P4CMDINSTR_P4CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P4CMDRA_P4CMDCLK_posedge : VitalTimingDataArrayType(14 downto 0);
      variable Tmkr_P4EN_P4CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P4WRDATA_P4CLK_posedge : VitalTimingDataArrayType(31 downto 0);
      variable Tmkr_P4WRMASK_P4CLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_P5ARBEN_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_P5CMDBA_P5CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P5CMDBL_P5CMDCLK_posedge : VitalTimingDataArrayType(5 downto 0);
      variable Tmkr_P5CMDCA_P5CMDCLK_posedge : VitalTimingDataArrayType(11 downto 0);
      variable Tmkr_P5CMDEN_P5CMDCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P5CMDINSTR_P5CMDCLK_posedge : VitalTimingDataArrayType(2 downto 0);
      variable Tmkr_P5CMDRA_P5CMDCLK_posedge : VitalTimingDataArrayType(14 downto 0);
      variable Tmkr_P5EN_P5CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_P5WRDATA_P5CLK_posedge : VitalTimingDataArrayType(31 downto 0);
      variable Tmkr_P5WRMASK_P5CLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_PLLCE_PLLCLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_PLLLOCK_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_RECAL_PLLCLK_posedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_SELFREFRESHENTER_PLLCLK_negedge : VitalTimingDataArrayType(1 downto 0);
      variable Tmkr_UIADDR_UICLK_posedge : VitalTimingDataArrayType(4 downto 0);
      variable Tmkr_UIADD_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIBROADCAST_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UICMDEN_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UICMDIN_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UICMD_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UICS_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIDONECAL_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIDQCOUNT_UICLK_posedge : VitalTimingDataArrayType(3 downto 0);
      variable Tmkr_UIDQLOWERDEC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIDQLOWERINC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIDQUPPERDEC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIDQUPPERINC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIDRPUPDATE_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UILDQSDEC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UILDQSINC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIREAD_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UISDI_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIUDQSDEC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Tmkr_UIUDQSINC_UICLK_posedge : VitalTimingDataType := VitalTimingDataInit;
      variable Pviol_PLLCLK : std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_IOIDRPSDI_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_P0ARBEN_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_P0CMDBA_P0CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P0CMDBL_P0CMDCLK_posedge : std_logic_vector(5 downto 0) := (others => '0');
      variable Tviol_P0CMDCA_P0CMDCLK_posedge : std_logic_vector(11 downto 0) := (others => '0');
      variable Tviol_P0CMDEN_P0CMDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P0CMDINSTR_P0CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P0CMDRA_P0CMDCLK_posedge : std_logic_vector(14 downto 0) := (others => '0');
      variable Tviol_P0RDEN_P0RDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P0RWRMASK_P0WRCLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_P0WRDATA_P0WRCLK_posedge : std_logic_vector(31 downto 0) := (others => '0');
      variable Tviol_P0WREN_P0WRCLK_posedge :  std_ulogic := '0';
      variable Tviol_P1ARBEN_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_P1CMDBA_P1CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P1CMDBL_P1CMDCLK_posedge : std_logic_vector(5 downto 0) := (others => '0');
      variable Tviol_P1CMDCA_P1CMDCLK_posedge : std_logic_vector(11 downto 0) := (others => '0');
      variable Tviol_P1CMDEN_P1CMDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P1CMDINSTR_P1CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P1CMDRA_P1CMDCLK_posedge : std_logic_vector(14 downto 0) := (others => '0');
      variable Tviol_P1RDEN_P1RDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P1RWRMASK_P1WRCLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_P1WRDATA_P1WRCLK_posedge : std_logic_vector(31 downto 0) := (others => '0');
      variable Tviol_P1WREN_P1WRCLK_posedge :  std_ulogic := '0';
      variable Tviol_P2ARBEN_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_P2CMDBA_P2CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P2CMDBL_P2CMDCLK_posedge : std_logic_vector(5 downto 0) := (others => '0');
      variable Tviol_P2CMDCA_P2CMDCLK_posedge : std_logic_vector(11 downto 0) := (others => '0');
      variable Tviol_P2CMDEN_P2CMDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P2CMDINSTR_P2CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P2CMDRA_P2CMDCLK_posedge : std_logic_vector(14 downto 0) := (others => '0');
      variable Tviol_P2EN_P2CLK_posedge :  std_ulogic := '0';
      variable Tviol_P2WRDATA_P2CLK_posedge : std_logic_vector(31 downto 0) := (others => '0');
      variable Tviol_P2WRMASK_P2CLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_P3ARBEN_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_P3CMDBA_P3CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P3CMDBL_P3CMDCLK_posedge : std_logic_vector(5 downto 0) := (others => '0');
      variable Tviol_P3CMDCA_P3CMDCLK_posedge : std_logic_vector(11 downto 0) := (others => '0');
      variable Tviol_P3CMDEN_P3CMDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P3CMDINSTR_P3CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P3CMDRA_P3CMDCLK_posedge : std_logic_vector(14 downto 0) := (others => '0');
      variable Tviol_P3EN_P3CLK_posedge :  std_ulogic := '0';
      variable Tviol_P3WRDATA_P3CLK_posedge : std_logic_vector(31 downto 0) := (others => '0');
      variable Tviol_P3WRMASK_P3CLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_P4ARBEN_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_P4CMDBA_P4CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P4CMDBL_P4CMDCLK_posedge : std_logic_vector(5 downto 0) := (others => '0');
      variable Tviol_P4CMDCA_P4CMDCLK_posedge : std_logic_vector(11 downto 0) := (others => '0');
      variable Tviol_P4CMDEN_P4CMDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P4CMDINSTR_P4CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P4CMDRA_P4CMDCLK_posedge : std_logic_vector(14 downto 0) := (others => '0');
      variable Tviol_P4EN_P4CLK_posedge :  std_ulogic := '0';
      variable Tviol_P4WRDATA_P4CLK_posedge : std_logic_vector(31 downto 0) := (others => '0');
      variable Tviol_P4WRMASK_P4CLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_P5ARBEN_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_P5CMDBA_P5CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P5CMDBL_P5CMDCLK_posedge : std_logic_vector(5 downto 0) := (others => '0');
      variable Tviol_P5CMDCA_P5CMDCLK_posedge : std_logic_vector(11 downto 0) := (others => '0');
      variable Tviol_P5CMDEN_P5CMDCLK_posedge :  std_ulogic := '0';
      variable Tviol_P5CMDINSTR_P5CMDCLK_posedge : std_logic_vector(2 downto 0) := (others => '0');
      variable Tviol_P5CMDRA_P5CMDCLK_posedge : std_logic_vector(14 downto 0) := (others => '0');
      variable Tviol_P5EN_P5CLK_posedge :  std_ulogic := '0';
      variable Tviol_P5WRDATA_P5CLK_posedge : std_logic_vector(31 downto 0) := (others => '0');
      variable Tviol_P5WRMASK_P5CLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_PLLCE_PLLCLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_PLLLOCK_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_RECAL_PLLCLK_posedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_SELFREFRESHENTER_PLLCLK_negedge :  std_logic_vector(1 downto 0) := (others => '0');
      variable Tviol_UIADDR_UICLK_posedge : std_logic_vector(4 downto 0) := (others => '0');
      variable Tviol_UIADD_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIBROADCAST_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UICMDEN_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UICMDIN_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UICMD_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UICS_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIDONECAL_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIDQCOUNT_UICLK_posedge : std_logic_vector(3 downto 0) := (others => '0');
      variable Tviol_UIDQLOWERDEC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIDQLOWERINC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIDQUPPERDEC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIDQUPPERINC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIDRPUPDATE_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UILDQSDEC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UILDQSINC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIREAD_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UISDI_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIUDQSDEC_UICLK_posedge :  std_ulogic := '0';
      variable Tviol_UIUDQSINC_UICLK_posedge :  std_ulogic := '0';
      variable DQIOWEN0_GlitchData : VitalGlitchDataType;
      variable DQSIOWEN90N_GlitchData : VitalGlitchDataType;
      variable DQSIOWEN90P_GlitchData : VitalGlitchDataType;
      variable IOIDRPADDR0_GlitchData : VitalGlitchDataType;
      variable IOIDRPADDR1_GlitchData : VitalGlitchDataType;
      variable IOIDRPADDR2_GlitchData : VitalGlitchDataType;
      variable IOIDRPADDR3_GlitchData : VitalGlitchDataType;
      variable IOIDRPADDR4_GlitchData : VitalGlitchDataType;
      variable IOIDRPADD_GlitchData : VitalGlitchDataType;
      variable IOIDRPBROADCAST_GlitchData : VitalGlitchDataType;
      variable IOIDRPCLK_GlitchData : VitalGlitchDataType;
      variable IOIDRPCS_GlitchData : VitalGlitchDataType;
      variable IOIDRPSDO_GlitchData : VitalGlitchDataType;
      variable IOIDRPUPDATE_GlitchData : VitalGlitchDataType;
      variable P0CMDEMPTY_GlitchData : VitalGlitchDataType;
      variable P0CMDFULL_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT0_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT1_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT2_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT3_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT4_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT5_GlitchData : VitalGlitchDataType;
      variable P0RDCOUNT6_GlitchData : VitalGlitchDataType;
      variable P0RDDATA0_GlitchData : VitalGlitchDataType;
      variable P0RDDATA10_GlitchData : VitalGlitchDataType;
      variable P0RDDATA11_GlitchData : VitalGlitchDataType;
      variable P0RDDATA12_GlitchData : VitalGlitchDataType;
      variable P0RDDATA13_GlitchData : VitalGlitchDataType;
      variable P0RDDATA14_GlitchData : VitalGlitchDataType;
      variable P0RDDATA15_GlitchData : VitalGlitchDataType;
      variable P0RDDATA16_GlitchData : VitalGlitchDataType;
      variable P0RDDATA17_GlitchData : VitalGlitchDataType;
      variable P0RDDATA18_GlitchData : VitalGlitchDataType;
      variable P0RDDATA19_GlitchData : VitalGlitchDataType;
      variable P0RDDATA1_GlitchData : VitalGlitchDataType;
      variable P0RDDATA20_GlitchData : VitalGlitchDataType;
      variable P0RDDATA21_GlitchData : VitalGlitchDataType;
      variable P0RDDATA22_GlitchData : VitalGlitchDataType;
      variable P0RDDATA23_GlitchData : VitalGlitchDataType;
      variable P0RDDATA24_GlitchData : VitalGlitchDataType;
      variable P0RDDATA25_GlitchData : VitalGlitchDataType;
      variable P0RDDATA26_GlitchData : VitalGlitchDataType;
      variable P0RDDATA27_GlitchData : VitalGlitchDataType;
      variable P0RDDATA28_GlitchData : VitalGlitchDataType;
      variable P0RDDATA29_GlitchData : VitalGlitchDataType;
      variable P0RDDATA2_GlitchData : VitalGlitchDataType;
      variable P0RDDATA30_GlitchData : VitalGlitchDataType;
      variable P0RDDATA31_GlitchData : VitalGlitchDataType;
      variable P0RDDATA3_GlitchData : VitalGlitchDataType;
      variable P0RDDATA4_GlitchData : VitalGlitchDataType;
      variable P0RDDATA5_GlitchData : VitalGlitchDataType;
      variable P0RDDATA6_GlitchData : VitalGlitchDataType;
      variable P0RDDATA7_GlitchData : VitalGlitchDataType;
      variable P0RDDATA8_GlitchData : VitalGlitchDataType;
      variable P0RDDATA9_GlitchData : VitalGlitchDataType;
      variable P0RDEMPTY_GlitchData : VitalGlitchDataType;
      variable P0RDERROR_GlitchData : VitalGlitchDataType;
      variable P0RDFULL_GlitchData : VitalGlitchDataType;
      variable P0RDOVERFLOW_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT0_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT1_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT2_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT3_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT4_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT5_GlitchData : VitalGlitchDataType;
      variable P0WRCOUNT6_GlitchData : VitalGlitchDataType;
      variable P0WREMPTY_GlitchData : VitalGlitchDataType;
      variable P0WRERROR_GlitchData : VitalGlitchDataType;
      variable P0WRFULL_GlitchData : VitalGlitchDataType;
      variable P0WRUNDERRUN_GlitchData : VitalGlitchDataType;
      variable P1CMDEMPTY_GlitchData : VitalGlitchDataType;
      variable P1CMDFULL_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT0_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT1_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT2_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT3_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT4_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT5_GlitchData : VitalGlitchDataType;
      variable P1RDCOUNT6_GlitchData : VitalGlitchDataType;
      variable P1RDDATA0_GlitchData : VitalGlitchDataType;
      variable P1RDDATA10_GlitchData : VitalGlitchDataType;
      variable P1RDDATA11_GlitchData : VitalGlitchDataType;
      variable P1RDDATA12_GlitchData : VitalGlitchDataType;
      variable P1RDDATA13_GlitchData : VitalGlitchDataType;
      variable P1RDDATA14_GlitchData : VitalGlitchDataType;
      variable P1RDDATA15_GlitchData : VitalGlitchDataType;
      variable P1RDDATA16_GlitchData : VitalGlitchDataType;
      variable P1RDDATA17_GlitchData : VitalGlitchDataType;
      variable P1RDDATA18_GlitchData : VitalGlitchDataType;
      variable P1RDDATA19_GlitchData : VitalGlitchDataType;
      variable P1RDDATA1_GlitchData : VitalGlitchDataType;
      variable P1RDDATA20_GlitchData : VitalGlitchDataType;
      variable P1RDDATA21_GlitchData : VitalGlitchDataType;
      variable P1RDDATA22_GlitchData : VitalGlitchDataType;
      variable P1RDDATA23_GlitchData : VitalGlitchDataType;
      variable P1RDDATA24_GlitchData : VitalGlitchDataType;
      variable P1RDDATA25_GlitchData : VitalGlitchDataType;
      variable P1RDDATA26_GlitchData : VitalGlitchDataType;
      variable P1RDDATA27_GlitchData : VitalGlitchDataType;
      variable P1RDDATA28_GlitchData : VitalGlitchDataType;
      variable P1RDDATA29_GlitchData : VitalGlitchDataType;
      variable P1RDDATA2_GlitchData : VitalGlitchDataType;
      variable P1RDDATA30_GlitchData : VitalGlitchDataType;
      variable P1RDDATA31_GlitchData : VitalGlitchDataType;
      variable P1RDDATA3_GlitchData : VitalGlitchDataType;
      variable P1RDDATA4_GlitchData : VitalGlitchDataType;
      variable P1RDDATA5_GlitchData : VitalGlitchDataType;
      variable P1RDDATA6_GlitchData : VitalGlitchDataType;
      variable P1RDDATA7_GlitchData : VitalGlitchDataType;
      variable P1RDDATA8_GlitchData : VitalGlitchDataType;
      variable P1RDDATA9_GlitchData : VitalGlitchDataType;
      variable P1RDEMPTY_GlitchData : VitalGlitchDataType;
      variable P1RDERROR_GlitchData : VitalGlitchDataType;
      variable P1RDFULL_GlitchData : VitalGlitchDataType;
      variable P1RDOVERFLOW_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT0_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT1_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT2_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT3_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT4_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT5_GlitchData : VitalGlitchDataType;
      variable P1WRCOUNT6_GlitchData : VitalGlitchDataType;
      variable P1WREMPTY_GlitchData : VitalGlitchDataType;
      variable P1WRERROR_GlitchData : VitalGlitchDataType;
      variable P1WRFULL_GlitchData : VitalGlitchDataType;
      variable P1WRUNDERRUN_GlitchData : VitalGlitchDataType;
      variable P2CMDEMPTY_GlitchData : VitalGlitchDataType;
      variable P2CMDFULL_GlitchData : VitalGlitchDataType;
      variable P2COUNT0_GlitchData : VitalGlitchDataType;
      variable P2COUNT1_GlitchData : VitalGlitchDataType;
      variable P2COUNT2_GlitchData : VitalGlitchDataType;
      variable P2COUNT3_GlitchData : VitalGlitchDataType;
      variable P2COUNT4_GlitchData : VitalGlitchDataType;
      variable P2COUNT5_GlitchData : VitalGlitchDataType;
      variable P2COUNT6_GlitchData : VitalGlitchDataType;
      variable P2EMPTY_GlitchData : VitalGlitchDataType;
      variable P2ERROR_GlitchData : VitalGlitchDataType;
      variable P2FULL_GlitchData : VitalGlitchDataType;
      variable P2RDDATA0_GlitchData : VitalGlitchDataType;
      variable P2RDDATA10_GlitchData : VitalGlitchDataType;
      variable P2RDDATA11_GlitchData : VitalGlitchDataType;
      variable P2RDDATA12_GlitchData : VitalGlitchDataType;
      variable P2RDDATA13_GlitchData : VitalGlitchDataType;
      variable P2RDDATA14_GlitchData : VitalGlitchDataType;
      variable P2RDDATA15_GlitchData : VitalGlitchDataType;
      variable P2RDDATA16_GlitchData : VitalGlitchDataType;
      variable P2RDDATA17_GlitchData : VitalGlitchDataType;
      variable P2RDDATA18_GlitchData : VitalGlitchDataType;
      variable P2RDDATA19_GlitchData : VitalGlitchDataType;
      variable P2RDDATA1_GlitchData : VitalGlitchDataType;
      variable P2RDDATA20_GlitchData : VitalGlitchDataType;
      variable P2RDDATA21_GlitchData : VitalGlitchDataType;
      variable P2RDDATA22_GlitchData : VitalGlitchDataType;
      variable P2RDDATA23_GlitchData : VitalGlitchDataType;
      variable P2RDDATA24_GlitchData : VitalGlitchDataType;
      variable P2RDDATA25_GlitchData : VitalGlitchDataType;
      variable P2RDDATA26_GlitchData : VitalGlitchDataType;
      variable P2RDDATA27_GlitchData : VitalGlitchDataType;
      variable P2RDDATA28_GlitchData : VitalGlitchDataType;
      variable P2RDDATA29_GlitchData : VitalGlitchDataType;
      variable P2RDDATA2_GlitchData : VitalGlitchDataType;
      variable P2RDDATA30_GlitchData : VitalGlitchDataType;
      variable P2RDDATA31_GlitchData : VitalGlitchDataType;
      variable P2RDDATA3_GlitchData : VitalGlitchDataType;
      variable P2RDDATA4_GlitchData : VitalGlitchDataType;
      variable P2RDDATA5_GlitchData : VitalGlitchDataType;
      variable P2RDDATA6_GlitchData : VitalGlitchDataType;
      variable P2RDDATA7_GlitchData : VitalGlitchDataType;
      variable P2RDDATA8_GlitchData : VitalGlitchDataType;
      variable P2RDDATA9_GlitchData : VitalGlitchDataType;
      variable P2RDOVERFLOW_GlitchData : VitalGlitchDataType;
      variable P2WRUNDERRUN_GlitchData : VitalGlitchDataType;
      variable P3CMDEMPTY_GlitchData : VitalGlitchDataType;
      variable P3CMDFULL_GlitchData : VitalGlitchDataType;
      variable P3COUNT0_GlitchData : VitalGlitchDataType;
      variable P3COUNT1_GlitchData : VitalGlitchDataType;
      variable P3COUNT2_GlitchData : VitalGlitchDataType;
      variable P3COUNT3_GlitchData : VitalGlitchDataType;
      variable P3COUNT4_GlitchData : VitalGlitchDataType;
      variable P3COUNT5_GlitchData : VitalGlitchDataType;
      variable P3COUNT6_GlitchData : VitalGlitchDataType;
      variable P3EMPTY_GlitchData : VitalGlitchDataType;
      variable P3ERROR_GlitchData : VitalGlitchDataType;
      variable P3FULL_GlitchData : VitalGlitchDataType;
      variable P3RDDATA0_GlitchData : VitalGlitchDataType;
      variable P3RDDATA10_GlitchData : VitalGlitchDataType;
      variable P3RDDATA11_GlitchData : VitalGlitchDataType;
      variable P3RDDATA12_GlitchData : VitalGlitchDataType;
      variable P3RDDATA13_GlitchData : VitalGlitchDataType;
      variable P3RDDATA14_GlitchData : VitalGlitchDataType;
      variable P3RDDATA15_GlitchData : VitalGlitchDataType;
      variable P3RDDATA16_GlitchData : VitalGlitchDataType;
      variable P3RDDATA17_GlitchData : VitalGlitchDataType;
      variable P3RDDATA18_GlitchData : VitalGlitchDataType;
      variable P3RDDATA19_GlitchData : VitalGlitchDataType;
      variable P3RDDATA1_GlitchData : VitalGlitchDataType;
      variable P3RDDATA20_GlitchData : VitalGlitchDataType;
      variable P3RDDATA21_GlitchData : VitalGlitchDataType;
      variable P3RDDATA22_GlitchData : VitalGlitchDataType;
      variable P3RDDATA23_GlitchData : VitalGlitchDataType;
      variable P3RDDATA24_GlitchData : VitalGlitchDataType;
      variable P3RDDATA25_GlitchData : VitalGlitchDataType;
      variable P3RDDATA26_GlitchData : VitalGlitchDataType;
      variable P3RDDATA27_GlitchData : VitalGlitchDataType;
      variable P3RDDATA28_GlitchData : VitalGlitchDataType;
      variable P3RDDATA29_GlitchData : VitalGlitchDataType;
      variable P3RDDATA2_GlitchData : VitalGlitchDataType;
      variable P3RDDATA30_GlitchData : VitalGlitchDataType;
      variable P3RDDATA31_GlitchData : VitalGlitchDataType;
      variable P3RDDATA3_GlitchData : VitalGlitchDataType;
      variable P3RDDATA4_GlitchData : VitalGlitchDataType;
      variable P3RDDATA5_GlitchData : VitalGlitchDataType;
      variable P3RDDATA6_GlitchData : VitalGlitchDataType;
      variable P3RDDATA7_GlitchData : VitalGlitchDataType;
      variable P3RDDATA8_GlitchData : VitalGlitchDataType;
      variable P3RDDATA9_GlitchData : VitalGlitchDataType;
      variable P3RDOVERFLOW_GlitchData : VitalGlitchDataType;
      variable P3WRUNDERRUN_GlitchData : VitalGlitchDataType;
      variable P4CMDEMPTY_GlitchData : VitalGlitchDataType;
      variable P4CMDFULL_GlitchData : VitalGlitchDataType;
      variable P4COUNT0_GlitchData : VitalGlitchDataType;
      variable P4COUNT1_GlitchData : VitalGlitchDataType;
      variable P4COUNT2_GlitchData : VitalGlitchDataType;
      variable P4COUNT3_GlitchData : VitalGlitchDataType;
      variable P4COUNT4_GlitchData : VitalGlitchDataType;
      variable P4COUNT5_GlitchData : VitalGlitchDataType;
      variable P4COUNT6_GlitchData : VitalGlitchDataType;
      variable P4EMPTY_GlitchData : VitalGlitchDataType;
      variable P4ERROR_GlitchData : VitalGlitchDataType;
      variable P4FULL_GlitchData : VitalGlitchDataType;
      variable P4RDDATA0_GlitchData : VitalGlitchDataType;
      variable P4RDDATA10_GlitchData : VitalGlitchDataType;
      variable P4RDDATA11_GlitchData : VitalGlitchDataType;
      variable P4RDDATA12_GlitchData : VitalGlitchDataType;
      variable P4RDDATA13_GlitchData : VitalGlitchDataType;
      variable P4RDDATA14_GlitchData : VitalGlitchDataType;
      variable P4RDDATA15_GlitchData : VitalGlitchDataType;
      variable P4RDDATA16_GlitchData : VitalGlitchDataType;
      variable P4RDDATA17_GlitchData : VitalGlitchDataType;
      variable P4RDDATA18_GlitchData : VitalGlitchDataType;
      variable P4RDDATA19_GlitchData : VitalGlitchDataType;
      variable P4RDDATA1_GlitchData : VitalGlitchDataType;
      variable P4RDDATA20_GlitchData : VitalGlitchDataType;
      variable P4RDDATA21_GlitchData : VitalGlitchDataType;
      variable P4RDDATA22_GlitchData : VitalGlitchDataType;
      variable P4RDDATA23_GlitchData : VitalGlitchDataType;
      variable P4RDDATA24_GlitchData : VitalGlitchDataType;
      variable P4RDDATA25_GlitchData : VitalGlitchDataType;
      variable P4RDDATA26_GlitchData : VitalGlitchDataType;
      variable P4RDDATA27_GlitchData : VitalGlitchDataType;
      variable P4RDDATA28_GlitchData : VitalGlitchDataType;
      variable P4RDDATA29_GlitchData : VitalGlitchDataType;
      variable P4RDDATA2_GlitchData : VitalGlitchDataType;
      variable P4RDDATA30_GlitchData : VitalGlitchDataType;
      variable P4RDDATA31_GlitchData : VitalGlitchDataType;
      variable P4RDDATA3_GlitchData : VitalGlitchDataType;
      variable P4RDDATA4_GlitchData : VitalGlitchDataType;
      variable P4RDDATA5_GlitchData : VitalGlitchDataType;
      variable P4RDDATA6_GlitchData : VitalGlitchDataType;
      variable P4RDDATA7_GlitchData : VitalGlitchDataType;
      variable P4RDDATA8_GlitchData : VitalGlitchDataType;
      variable P4RDDATA9_GlitchData : VitalGlitchDataType;
      variable P4RDOVERFLOW_GlitchData : VitalGlitchDataType;
      variable P4WRUNDERRUN_GlitchData : VitalGlitchDataType;
      variable P5CMDEMPTY_GlitchData : VitalGlitchDataType;
      variable P5CMDFULL_GlitchData : VitalGlitchDataType;
      variable P5COUNT0_GlitchData : VitalGlitchDataType;
      variable P5COUNT1_GlitchData : VitalGlitchDataType;
      variable P5COUNT2_GlitchData : VitalGlitchDataType;
      variable P5COUNT3_GlitchData : VitalGlitchDataType;
      variable P5COUNT4_GlitchData : VitalGlitchDataType;
      variable P5COUNT5_GlitchData : VitalGlitchDataType;
      variable P5COUNT6_GlitchData : VitalGlitchDataType;
      variable P5EMPTY_GlitchData : VitalGlitchDataType;
      variable P5ERROR_GlitchData : VitalGlitchDataType;
      variable P5FULL_GlitchData : VitalGlitchDataType;
      variable P5RDDATA0_GlitchData : VitalGlitchDataType;
      variable P5RDDATA10_GlitchData : VitalGlitchDataType;
      variable P5RDDATA11_GlitchData : VitalGlitchDataType;
      variable P5RDDATA12_GlitchData : VitalGlitchDataType;
      variable P5RDDATA13_GlitchData : VitalGlitchDataType;
      variable P5RDDATA14_GlitchData : VitalGlitchDataType;
      variable P5RDDATA15_GlitchData : VitalGlitchDataType;
      variable P5RDDATA16_GlitchData : VitalGlitchDataType;
      variable P5RDDATA17_GlitchData : VitalGlitchDataType;
      variable P5RDDATA18_GlitchData : VitalGlitchDataType;
      variable P5RDDATA19_GlitchData : VitalGlitchDataType;
      variable P5RDDATA1_GlitchData : VitalGlitchDataType;
      variable P5RDDATA20_GlitchData : VitalGlitchDataType;
      variable P5RDDATA21_GlitchData : VitalGlitchDataType;
      variable P5RDDATA22_GlitchData : VitalGlitchDataType;
      variable P5RDDATA23_GlitchData : VitalGlitchDataType;
      variable P5RDDATA24_GlitchData : VitalGlitchDataType;
      variable P5RDDATA25_GlitchData : VitalGlitchDataType;
      variable P5RDDATA26_GlitchData : VitalGlitchDataType;
      variable P5RDDATA27_GlitchData : VitalGlitchDataType;
      variable P5RDDATA28_GlitchData : VitalGlitchDataType;
      variable P5RDDATA29_GlitchData : VitalGlitchDataType;
      variable P5RDDATA2_GlitchData : VitalGlitchDataType;
      variable P5RDDATA30_GlitchData : VitalGlitchDataType;
      variable P5RDDATA31_GlitchData : VitalGlitchDataType;
      variable P5RDDATA3_GlitchData : VitalGlitchDataType;
      variable P5RDDATA4_GlitchData : VitalGlitchDataType;
      variable P5RDDATA5_GlitchData : VitalGlitchDataType;
      variable P5RDDATA6_GlitchData : VitalGlitchDataType;
      variable P5RDDATA7_GlitchData : VitalGlitchDataType;
      variable P5RDDATA8_GlitchData : VitalGlitchDataType;
      variable P5RDDATA9_GlitchData : VitalGlitchDataType;
      variable P5RDOVERFLOW_GlitchData : VitalGlitchDataType;
      variable P5WRUNDERRUN_GlitchData : VitalGlitchDataType;
      variable SELFREFRESHMODE_GlitchData : VitalGlitchDataType;
      variable UOCALSTART_GlitchData : VitalGlitchDataType;
      variable UOCMDREADYIN_GlitchData : VitalGlitchDataType;
      variable UODATA0_GlitchData : VitalGlitchDataType;
      variable UODATA1_GlitchData : VitalGlitchDataType;
      variable UODATA2_GlitchData : VitalGlitchDataType;
      variable UODATA3_GlitchData : VitalGlitchDataType;
      variable UODATA4_GlitchData : VitalGlitchDataType;
      variable UODATA5_GlitchData : VitalGlitchDataType;
      variable UODATA6_GlitchData : VitalGlitchDataType;
      variable UODATA7_GlitchData : VitalGlitchDataType;
      variable UODATAVALID_GlitchData : VitalGlitchDataType;
      variable UODONECAL_GlitchData : VitalGlitchDataType;
      variable UOREFRSHFLAG_GlitchData : VitalGlitchDataType;
      variable UOSDO_GlitchData : VitalGlitchDataType;
      variable Pviol_P0CMDCLK : STD_ULOGIC := '0';
      variable Pviol_P0RDCLK : STD_ULOGIC := '0';
      variable Pviol_P0WRCLK : STD_ULOGIC := '0';
      variable Pviol_P1CMDCLK : STD_ULOGIC := '0';
      variable Pviol_P1RDCLK : STD_ULOGIC := '0';
      variable Pviol_P1WRCLK : STD_ULOGIC := '0';
      variable Pviol_P2CLK : STD_ULOGIC := '0';
      variable Pviol_P2CMDCLK : STD_ULOGIC := '0';
      variable Pviol_P3CLK : STD_ULOGIC := '0';
      variable Pviol_P3CMDCLK : STD_ULOGIC := '0';
      variable Pviol_P4CLK : STD_ULOGIC := '0';
      variable Pviol_P4CMDCLK : STD_ULOGIC := '0';
      variable Pviol_P5CLK : STD_ULOGIC := '0';
      variable Pviol_P5CMDCLK : STD_ULOGIC := '0';
      variable Pviol_SYSRST : STD_ULOGIC := '0';
      variable Pviol_UICLK : STD_ULOGIC := '0';
      variable PInfo_P0CMDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P0RDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P0WRCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P1CMDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P1RDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P1WRCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P2CLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P2CMDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P3CLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P3CMDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P4CLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P4CMDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P5CLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_P5CMDCLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_SYSRST : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_UICLK : VitalPeriodDataType := VitalPeriodDataInit;
      variable PInfo_PLLCLK : VitalPeriodDataType := VitalPeriodDataInit;

      begin

      if (TimingChecksOn) then
        VitalSetupHoldCheck
        (
          Violation => Tviol_IOIDRPSDI_UICLK_posedge,
          TimingData => Tmkr_IOIDRPSDI_UICLK_posedge,
          TestSignal => IOIDRPSDI_UICLK_dly,
          TestSignalName => "IOIDRPSDI",
          TestDelay => tisd_IOIDRPSDI_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_IOIDRPSDI_UICLK_posedge_posedge,
          HoldHigh => thold_IOIDRPSDI_UICLK_posedge_posedge,
          SetupLow => tsetup_IOIDRPSDI_UICLK_negedge_posedge,
          HoldLow => thold_IOIDRPSDI_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
       VitalSetupHoldCheck
        (
          Violation => Tviol_P0ARBEN_PLLCLK_posedge(0),
          TimingData => Tmkr_P0ARBEN_PLLCLK_posedge(0),
          TestSignal => P0ARBEN_PLLCLK_dly(0),
          TestSignalName => "P0ARBEN",
          TestDelay => tisd_P0ARBEN_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_P0ARBEN_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_P0ARBEN_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_P0ARBEN_PLLCLK_negedge_posedge(0),
          HoldLow => thold_P0ARBEN_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0ARBEN_PLLCLK_posedge(1),
          TimingData => Tmkr_P0ARBEN_PLLCLK_posedge(1),
          TestSignal => P0ARBEN_PLLCLK_dly(1),
          TestSignalName => "P0ARBEN",
          TestDelay => tisd_P0ARBEN_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_P0ARBEN_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_P0ARBEN_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_P0ARBEN_PLLCLK_negedge_posedge(1),
          HoldLow => thold_P0ARBEN_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
       
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBA_P0CMDCLK_posedge(0),
          TimingData => Tmkr_P0CMDBA_P0CMDCLK_posedge(0),
          TestSignal => P0CMDBA_P0CMDCLK_dly(0),
          TestSignalName => "P0CMDBA(0)",
          TestDelay => tisd_P0CMDBA_P0CMDCLK(0),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBA_P0CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P0CMDBA_P0CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P0CMDBA_P0CMDCLK_negedge_posedge(0),
          HoldLow => thold_P0CMDBA_P0CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBA_P0CMDCLK_posedge(1),
          TimingData => Tmkr_P0CMDBA_P0CMDCLK_posedge(1),
          TestSignal => P0CMDBA_P0CMDCLK_dly(1),
          TestSignalName => "P0CMDBA(1)",
          TestDelay => tisd_P0CMDBA_P0CMDCLK(1),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBA_P0CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P0CMDBA_P0CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P0CMDBA_P0CMDCLK_negedge_posedge(1),
          HoldLow => thold_P0CMDBA_P0CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBA_P0CMDCLK_posedge(2),
          TimingData => Tmkr_P0CMDBA_P0CMDCLK_posedge(2),
          TestSignal => P0CMDBA_P0CMDCLK_dly(2),
          TestSignalName => "P0CMDBA(2)",
          TestDelay => tisd_P0CMDBA_P0CMDCLK(2),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBA_P0CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P0CMDBA_P0CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P0CMDBA_P0CMDCLK_negedge_posedge(2),
          HoldLow => thold_P0CMDBA_P0CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBL_P0CMDCLK_posedge(0),
          TimingData => Tmkr_P0CMDBL_P0CMDCLK_posedge(0),
          TestSignal => P0CMDBL_P0CMDCLK_dly(0),
          TestSignalName => "P0CMDBL(0)",
          TestDelay => tisd_P0CMDBL_P0CMDCLK(0),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBL_P0CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P0CMDBL_P0CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P0CMDBL_P0CMDCLK_negedge_posedge(0),
          HoldLow => thold_P0CMDBL_P0CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBL_P0CMDCLK_posedge(1),
          TimingData => Tmkr_P0CMDBL_P0CMDCLK_posedge(1),
          TestSignal => P0CMDBL_P0CMDCLK_dly(1),
          TestSignalName => "P0CMDBL(1)",
          TestDelay => tisd_P0CMDBL_P0CMDCLK(1),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBL_P0CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P0CMDBL_P0CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P0CMDBL_P0CMDCLK_negedge_posedge(1),
          HoldLow => thold_P0CMDBL_P0CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBL_P0CMDCLK_posedge(2),
          TimingData => Tmkr_P0CMDBL_P0CMDCLK_posedge(2),
          TestSignal => P0CMDBL_P0CMDCLK_dly(2),
          TestSignalName => "P0CMDBL(2)",
          TestDelay => tisd_P0CMDBL_P0CMDCLK(2),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBL_P0CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P0CMDBL_P0CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P0CMDBL_P0CMDCLK_negedge_posedge(2),
          HoldLow => thold_P0CMDBL_P0CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBL_P0CMDCLK_posedge(3),
          TimingData => Tmkr_P0CMDBL_P0CMDCLK_posedge(3),
          TestSignal => P0CMDBL_P0CMDCLK_dly(3),
          TestSignalName => "P0CMDBL(3)",
          TestDelay => tisd_P0CMDBL_P0CMDCLK(3),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBL_P0CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P0CMDBL_P0CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P0CMDBL_P0CMDCLK_negedge_posedge(3),
          HoldLow => thold_P0CMDBL_P0CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBL_P0CMDCLK_posedge(4),
          TimingData => Tmkr_P0CMDBL_P0CMDCLK_posedge(4),
          TestSignal => P0CMDBL_P0CMDCLK_dly(4),
          TestSignalName => "P0CMDBL(4)",
          TestDelay => tisd_P0CMDBL_P0CMDCLK(4),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBL_P0CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P0CMDBL_P0CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P0CMDBL_P0CMDCLK_negedge_posedge(4),
          HoldLow => thold_P0CMDBL_P0CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDBL_P0CMDCLK_posedge(5),
          TimingData => Tmkr_P0CMDBL_P0CMDCLK_posedge(5),
          TestSignal => P0CMDBL_P0CMDCLK_dly(5),
          TestSignalName => "P0CMDBL(5)",
          TestDelay => tisd_P0CMDBL_P0CMDCLK(5),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDBL_P0CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P0CMDBL_P0CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P0CMDBL_P0CMDCLK_negedge_posedge(5),
          HoldLow => thold_P0CMDBL_P0CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(0),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(0),
          TestSignal => P0CMDCA_P0CMDCLK_dly(0),
          TestSignalName => "P0CMDCA(0)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(0),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(0),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(1),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(1),
          TestSignal => P0CMDCA_P0CMDCLK_dly(1),
          TestSignalName => "P0CMDCA(1)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(1),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(1),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(10),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(10),
          TestSignal => P0CMDCA_P0CMDCLK_dly(10),
          TestSignalName => "P0CMDCA(10)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(10),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(10),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(11),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(11),
          TestSignal => P0CMDCA_P0CMDCLK_dly(11),
          TestSignalName => "P0CMDCA(11)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(11),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(11),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(2),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(2),
          TestSignal => P0CMDCA_P0CMDCLK_dly(2),
          TestSignalName => "P0CMDCA(2)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(2),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(2),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(3),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(3),
          TestSignal => P0CMDCA_P0CMDCLK_dly(3),
          TestSignalName => "P0CMDCA(3)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(3),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(3),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(4),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(4),
          TestSignal => P0CMDCA_P0CMDCLK_dly(4),
          TestSignalName => "P0CMDCA(4)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(4),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(4),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(5),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(5),
          TestSignal => P0CMDCA_P0CMDCLK_dly(5),
          TestSignalName => "P0CMDCA(5)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(5),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(5),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(6),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(6),
          TestSignal => P0CMDCA_P0CMDCLK_dly(6),
          TestSignalName => "P0CMDCA(6)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(6),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(6),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(7),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(7),
          TestSignal => P0CMDCA_P0CMDCLK_dly(7),
          TestSignalName => "P0CMDCA(7)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(7),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(7),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(8),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(8),
          TestSignal => P0CMDCA_P0CMDCLK_dly(8),
          TestSignalName => "P0CMDCA(8)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(8),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(8),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDCA_P0CMDCLK_posedge(9),
          TimingData => Tmkr_P0CMDCA_P0CMDCLK_posedge(9),
          TestSignal => P0CMDCA_P0CMDCLK_dly(9),
          TestSignalName => "P0CMDCA(9)",
          TestDelay => tisd_P0CMDCA_P0CMDCLK(9),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDCA_P0CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P0CMDCA_P0CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P0CMDCA_P0CMDCLK_negedge_posedge(9),
          HoldLow => thold_P0CMDCA_P0CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDEN_P0CMDCLK_posedge,
          TimingData => Tmkr_P0CMDEN_P0CMDCLK_posedge,
          TestSignal => P0CMDEN_P0CMDCLK_dly,
          TestSignalName => "P0CMDEN",
          TestDelay => tisd_P0CMDEN_P0CMDCLK,
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDEN_P0CMDCLK_posedge_posedge,
          HoldHigh => thold_P0CMDEN_P0CMDCLK_posedge_posedge,
          SetupLow => tsetup_P0CMDEN_P0CMDCLK_negedge_posedge,
          HoldLow => thold_P0CMDEN_P0CMDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDINSTR_P0CMDCLK_posedge(0),
          TimingData => Tmkr_P0CMDINSTR_P0CMDCLK_posedge(0),
          TestSignal => P0CMDINSTR_P0CMDCLK_dly(0),
          TestSignalName => "P0CMDINSTR(0)",
          TestDelay => tisd_P0CMDINSTR_P0CMDCLK(0),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDINSTR_P0CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P0CMDINSTR_P0CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P0CMDINSTR_P0CMDCLK_negedge_posedge(0),
          HoldLow => thold_P0CMDINSTR_P0CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDINSTR_P0CMDCLK_posedge(1),
          TimingData => Tmkr_P0CMDINSTR_P0CMDCLK_posedge(1),
          TestSignal => P0CMDINSTR_P0CMDCLK_dly(1),
          TestSignalName => "P0CMDINSTR(1)",
          TestDelay => tisd_P0CMDINSTR_P0CMDCLK(1),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDINSTR_P0CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P0CMDINSTR_P0CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P0CMDINSTR_P0CMDCLK_negedge_posedge(1),
          HoldLow => thold_P0CMDINSTR_P0CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDINSTR_P0CMDCLK_posedge(2),
          TimingData => Tmkr_P0CMDINSTR_P0CMDCLK_posedge(2),
          TestSignal => P0CMDINSTR_P0CMDCLK_dly(2),
          TestSignalName => "P0CMDINSTR(2)",
          TestDelay => tisd_P0CMDINSTR_P0CMDCLK(2),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDINSTR_P0CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P0CMDINSTR_P0CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P0CMDINSTR_P0CMDCLK_negedge_posedge(2),
          HoldLow => thold_P0CMDINSTR_P0CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(0),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(0),
          TestSignal => P0CMDRA_P0CMDCLK_dly(0),
          TestSignalName => "P0CMDRA(0)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(0),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(0),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(1),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(1),
          TestSignal => P0CMDRA_P0CMDCLK_dly(1),
          TestSignalName => "P0CMDRA(1)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(1),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(1),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(10),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(10),
          TestSignal => P0CMDRA_P0CMDCLK_dly(10),
          TestSignalName => "P0CMDRA(10)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(10),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(10),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(11),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(11),
          TestSignal => P0CMDRA_P0CMDCLK_dly(11),
          TestSignalName => "P0CMDRA(11)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(11),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(11),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(12),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(12),
          TestSignal => P0CMDRA_P0CMDCLK_dly(12),
          TestSignalName => "P0CMDRA(12)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(12),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(12),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(12),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(12),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(13),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(13),
          TestSignal => P0CMDRA_P0CMDCLK_dly(13),
          TestSignalName => "P0CMDRA(13)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(13),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(13),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(13),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(13),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(14),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(14),
          TestSignal => P0CMDRA_P0CMDCLK_dly(14),
          TestSignalName => "P0CMDRA(14)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(14),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(14),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(14),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(14),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(2),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(2),
          TestSignal => P0CMDRA_P0CMDCLK_dly(2),
          TestSignalName => "P0CMDRA(2)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(2),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(2),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(3),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(3),
          TestSignal => P0CMDRA_P0CMDCLK_dly(3),
          TestSignalName => "P0CMDRA(3)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(3),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(3),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(4),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(4),
          TestSignal => P0CMDRA_P0CMDCLK_dly(4),
          TestSignalName => "P0CMDRA(4)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(4),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(4),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(5),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(5),
          TestSignal => P0CMDRA_P0CMDCLK_dly(5),
          TestSignalName => "P0CMDRA(5)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(5),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(5),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(6),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(6),
          TestSignal => P0CMDRA_P0CMDCLK_dly(6),
          TestSignalName => "P0CMDRA(6)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(6),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(6),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(7),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(7),
          TestSignal => P0CMDRA_P0CMDCLK_dly(7),
          TestSignalName => "P0CMDRA(7)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(7),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(7),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(8),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(8),
          TestSignal => P0CMDRA_P0CMDCLK_dly(8),
          TestSignalName => "P0CMDRA(8)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(8),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(8),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0CMDRA_P0CMDCLK_posedge(9),
          TimingData => Tmkr_P0CMDRA_P0CMDCLK_posedge(9),
          TestSignal => P0CMDRA_P0CMDCLK_dly(9),
          TestSignalName => "P0CMDRA(9)",
          TestDelay => tisd_P0CMDRA_P0CMDCLK(9),
          RefSignal => P0CMDCLK_dly,
          RefSignalName => "P0CMDCLK",
          RefDelay => ticd_P0CMDCLK,
          SetupHigh => tsetup_P0CMDRA_P0CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P0CMDRA_P0CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P0CMDRA_P0CMDCLK_negedge_posedge(9),
          HoldLow => thold_P0CMDRA_P0CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0RDEN_P0RDCLK_posedge,
          TimingData => Tmkr_P0RDEN_P0RDCLK_posedge,
          TestSignal => P0RDEN_P0RDCLK_dly,
          TestSignalName => "P0RDEN",
          TestDelay => tisd_P0RDEN_P0RDCLK,
          RefSignal => P0RDCLK_dly,
          RefSignalName => "P0RDCLK",
          RefDelay => ticd_P0RDCLK,
          SetupHigh => tsetup_P0RDEN_P0RDCLK_posedge_posedge,
          HoldHigh => thold_P0RDEN_P0RDCLK_posedge_posedge,
          SetupLow => tsetup_P0RDEN_P0RDCLK_negedge_posedge,
          HoldLow => thold_P0RDEN_P0RDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0RWRMASK_P0WRCLK_posedge(0),
          TimingData => Tmkr_P0RWRMASK_P0WRCLK_posedge(0),
          TestSignal => P0RWRMASK_P0WRCLK_dly(0),
          TestSignalName => "P0RWRMASK(0)",
          TestDelay => tisd_P0RWRMASK_P0WRCLK(0),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0RWRMASK_P0WRCLK_posedge_posedge(0),
          HoldHigh => thold_P0RWRMASK_P0WRCLK_posedge_posedge(0),
          SetupLow => tsetup_P0RWRMASK_P0WRCLK_negedge_posedge(0),
          HoldLow => thold_P0RWRMASK_P0WRCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0RWRMASK_P0WRCLK_posedge(1),
          TimingData => Tmkr_P0RWRMASK_P0WRCLK_posedge(1),
          TestSignal => P0RWRMASK_P0WRCLK_dly(1),
          TestSignalName => "P0RWRMASK(1)",
          TestDelay => tisd_P0RWRMASK_P0WRCLK(1),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0RWRMASK_P0WRCLK_posedge_posedge(1),
          HoldHigh => thold_P0RWRMASK_P0WRCLK_posedge_posedge(1),
          SetupLow => tsetup_P0RWRMASK_P0WRCLK_negedge_posedge(1),
          HoldLow => thold_P0RWRMASK_P0WRCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0RWRMASK_P0WRCLK_posedge(2),
          TimingData => Tmkr_P0RWRMASK_P0WRCLK_posedge(2),
          TestSignal => P0RWRMASK_P0WRCLK_dly(2),
          TestSignalName => "P0RWRMASK(2)",
          TestDelay => tisd_P0RWRMASK_P0WRCLK(2),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0RWRMASK_P0WRCLK_posedge_posedge(2),
          HoldHigh => thold_P0RWRMASK_P0WRCLK_posedge_posedge(2),
          SetupLow => tsetup_P0RWRMASK_P0WRCLK_negedge_posedge(2),
          HoldLow => thold_P0RWRMASK_P0WRCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0RWRMASK_P0WRCLK_posedge(3),
          TimingData => Tmkr_P0RWRMASK_P0WRCLK_posedge(3),
          TestSignal => P0RWRMASK_P0WRCLK_dly(3),
          TestSignalName => "P0RWRMASK(3)",
          TestDelay => tisd_P0RWRMASK_P0WRCLK(3),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0RWRMASK_P0WRCLK_posedge_posedge(3),
          HoldHigh => thold_P0RWRMASK_P0WRCLK_posedge_posedge(3),
          SetupLow => tsetup_P0RWRMASK_P0WRCLK_negedge_posedge(3),
          HoldLow => thold_P0RWRMASK_P0WRCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(0),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(0),
          TestSignal => P0WRDATA_P0WRCLK_dly(0),
          TestSignalName => "P0WRDATA(0)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(0),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(0),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(0),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(0),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(1),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(1),
          TestSignal => P0WRDATA_P0WRCLK_dly(1),
          TestSignalName => "P0WRDATA(1)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(1),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(1),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(1),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(1),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(10),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(10),
          TestSignal => P0WRDATA_P0WRCLK_dly(10),
          TestSignalName => "P0WRDATA(10)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(10),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(10),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(10),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(10),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(11),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(11),
          TestSignal => P0WRDATA_P0WRCLK_dly(11),
          TestSignalName => "P0WRDATA(11)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(11),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(11),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(11),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(11),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(12),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(12),
          TestSignal => P0WRDATA_P0WRCLK_dly(12),
          TestSignalName => "P0WRDATA(12)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(12),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(12),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(12),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(12),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(13),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(13),
          TestSignal => P0WRDATA_P0WRCLK_dly(13),
          TestSignalName => "P0WRDATA(13)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(13),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(13),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(13),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(13),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(14),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(14),
          TestSignal => P0WRDATA_P0WRCLK_dly(14),
          TestSignalName => "P0WRDATA(14)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(14),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(14),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(14),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(14),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(15),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(15),
          TestSignal => P0WRDATA_P0WRCLK_dly(15),
          TestSignalName => "P0WRDATA(15)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(15),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(15),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(15),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(15),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(15),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(16),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(16),
          TestSignal => P0WRDATA_P0WRCLK_dly(16),
          TestSignalName => "P0WRDATA(16)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(16),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(16),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(16),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(16),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(16),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(17),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(17),
          TestSignal => P0WRDATA_P0WRCLK_dly(17),
          TestSignalName => "P0WRDATA(17)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(17),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(17),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(17),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(17),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(17),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(18),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(18),
          TestSignal => P0WRDATA_P0WRCLK_dly(18),
          TestSignalName => "P0WRDATA(18)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(18),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(18),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(18),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(18),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(18),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(19),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(19),
          TestSignal => P0WRDATA_P0WRCLK_dly(19),
          TestSignalName => "P0WRDATA(19)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(19),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(19),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(19),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(19),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(19),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(2),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(2),
          TestSignal => P0WRDATA_P0WRCLK_dly(2),
          TestSignalName => "P0WRDATA(2)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(2),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(2),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(2),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(2),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(20),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(20),
          TestSignal => P0WRDATA_P0WRCLK_dly(20),
          TestSignalName => "P0WRDATA(20)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(20),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(20),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(20),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(20),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(20),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(21),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(21),
          TestSignal => P0WRDATA_P0WRCLK_dly(21),
          TestSignalName => "P0WRDATA(21)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(21),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(21),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(21),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(21),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(21),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(22),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(22),
          TestSignal => P0WRDATA_P0WRCLK_dly(22),
          TestSignalName => "P0WRDATA(22)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(22),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(22),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(22),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(22),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(22),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(23),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(23),
          TestSignal => P0WRDATA_P0WRCLK_dly(23),
          TestSignalName => "P0WRDATA(23)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(23),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(23),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(23),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(23),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(23),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(24),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(24),
          TestSignal => P0WRDATA_P0WRCLK_dly(24),
          TestSignalName => "P0WRDATA(24)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(24),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(24),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(24),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(24),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(24),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(25),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(25),
          TestSignal => P0WRDATA_P0WRCLK_dly(25),
          TestSignalName => "P0WRDATA(25)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(25),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(25),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(25),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(25),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(25),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(26),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(26),
          TestSignal => P0WRDATA_P0WRCLK_dly(26),
          TestSignalName => "P0WRDATA(26)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(26),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(26),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(26),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(26),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(26),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(27),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(27),
          TestSignal => P0WRDATA_P0WRCLK_dly(27),
          TestSignalName => "P0WRDATA(27)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(27),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(27),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(27),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(27),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(27),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(28),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(28),
          TestSignal => P0WRDATA_P0WRCLK_dly(28),
          TestSignalName => "P0WRDATA(28)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(28),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(28),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(28),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(28),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(28),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(29),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(29),
          TestSignal => P0WRDATA_P0WRCLK_dly(29),
          TestSignalName => "P0WRDATA(29)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(29),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(29),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(29),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(29),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(29),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(3),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(3),
          TestSignal => P0WRDATA_P0WRCLK_dly(3),
          TestSignalName => "P0WRDATA(3)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(3),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(3),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(3),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(3),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(30),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(30),
          TestSignal => P0WRDATA_P0WRCLK_dly(30),
          TestSignalName => "P0WRDATA(30)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(30),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(30),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(30),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(30),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(30),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(31),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(31),
          TestSignal => P0WRDATA_P0WRCLK_dly(31),
          TestSignalName => "P0WRDATA(31)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(31),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(31),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(31),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(31),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(31),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(4),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(4),
          TestSignal => P0WRDATA_P0WRCLK_dly(4),
          TestSignalName => "P0WRDATA(4)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(4),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(4),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(4),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(4),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(5),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(5),
          TestSignal => P0WRDATA_P0WRCLK_dly(5),
          TestSignalName => "P0WRDATA(5)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(5),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(5),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(5),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(5),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(6),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(6),
          TestSignal => P0WRDATA_P0WRCLK_dly(6),
          TestSignalName => "P0WRDATA(6)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(6),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(6),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(6),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(6),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(7),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(7),
          TestSignal => P0WRDATA_P0WRCLK_dly(7),
          TestSignalName => "P0WRDATA(7)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(7),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(7),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(7),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(7),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(8),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(8),
          TestSignal => P0WRDATA_P0WRCLK_dly(8),
          TestSignalName => "P0WRDATA(8)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(8),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(8),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(8),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(8),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WRDATA_P0WRCLK_posedge(9),
          TimingData => Tmkr_P0WRDATA_P0WRCLK_posedge(9),
          TestSignal => P0WRDATA_P0WRCLK_dly(9),
          TestSignalName => "P0WRDATA(9)",
          TestDelay => tisd_P0WRDATA_P0WRCLK(9),
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WRDATA_P0WRCLK_posedge_posedge(9),
          HoldHigh => thold_P0WRDATA_P0WRCLK_posedge_posedge(9),
          SetupLow => tsetup_P0WRDATA_P0WRCLK_negedge_posedge(9),
          HoldLow => thold_P0WRDATA_P0WRCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P0WREN_P0WRCLK_posedge,
          TimingData => Tmkr_P0WREN_P0WRCLK_posedge,
          TestSignal => P0WREN_P0WRCLK_dly,
          TestSignalName => "P0WREN",
          TestDelay => tisd_P0WREN_P0WRCLK,
          RefSignal => P0WRCLK_dly,
          RefSignalName => "P0WRCLK",
          RefDelay => ticd_P0WRCLK,
          SetupHigh => tsetup_P0WREN_P0WRCLK_posedge_posedge,
          HoldHigh => thold_P0WREN_P0WRCLK_posedge_posedge,
          SetupLow => tsetup_P0WREN_P0WRCLK_negedge_posedge,
          HoldLow => thold_P0WREN_P0WRCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
       VitalSetupHoldCheck
        (
          Violation => Tviol_P1ARBEN_PLLCLK_posedge(0),
          TimingData => Tmkr_P1ARBEN_PLLCLK_posedge(0),
          TestSignal => P1ARBEN_PLLCLK_dly(0),
          TestSignalName => "P1ARBEN",
          TestDelay => tisd_P1ARBEN_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_P1ARBEN_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_P1ARBEN_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_P1ARBEN_PLLCLK_negedge_posedge(0),
          HoldLow => thold_P1ARBEN_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1ARBEN_PLLCLK_posedge(1),
          TimingData => Tmkr_P1ARBEN_PLLCLK_posedge(1),
          TestSignal => P1ARBEN_PLLCLK_dly(1),
          TestSignalName => "P1ARBEN",
          TestDelay => tisd_P1ARBEN_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_P1ARBEN_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_P1ARBEN_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_P1ARBEN_PLLCLK_negedge_posedge(1),
          HoldLow => thold_P1ARBEN_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBA_P1CMDCLK_posedge(0),
          TimingData => Tmkr_P1CMDBA_P1CMDCLK_posedge(0),
          TestSignal => P1CMDBA_P1CMDCLK_dly(0),
          TestSignalName => "P1CMDBA(0)",
          TestDelay => tisd_P1CMDBA_P1CMDCLK(0),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBA_P1CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P1CMDBA_P1CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P1CMDBA_P1CMDCLK_negedge_posedge(0),
          HoldLow => thold_P1CMDBA_P1CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBA_P1CMDCLK_posedge(1),
          TimingData => Tmkr_P1CMDBA_P1CMDCLK_posedge(1),
          TestSignal => P1CMDBA_P1CMDCLK_dly(1),
          TestSignalName => "P1CMDBA(1)",
          TestDelay => tisd_P1CMDBA_P1CMDCLK(1),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBA_P1CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P1CMDBA_P1CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P1CMDBA_P1CMDCLK_negedge_posedge(1),
          HoldLow => thold_P1CMDBA_P1CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBA_P1CMDCLK_posedge(2),
          TimingData => Tmkr_P1CMDBA_P1CMDCLK_posedge(2),
          TestSignal => P1CMDBA_P1CMDCLK_dly(2),
          TestSignalName => "P1CMDBA(2)",
          TestDelay => tisd_P1CMDBA_P1CMDCLK(2),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBA_P1CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P1CMDBA_P1CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P1CMDBA_P1CMDCLK_negedge_posedge(2),
          HoldLow => thold_P1CMDBA_P1CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBL_P1CMDCLK_posedge(0),
          TimingData => Tmkr_P1CMDBL_P1CMDCLK_posedge(0),
          TestSignal => P1CMDBL_P1CMDCLK_dly(0),
          TestSignalName => "P1CMDBL(0)",
          TestDelay => tisd_P1CMDBL_P1CMDCLK(0),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBL_P1CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P1CMDBL_P1CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P1CMDBL_P1CMDCLK_negedge_posedge(0),
          HoldLow => thold_P1CMDBL_P1CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBL_P1CMDCLK_posedge(1),
          TimingData => Tmkr_P1CMDBL_P1CMDCLK_posedge(1),
          TestSignal => P1CMDBL_P1CMDCLK_dly(1),
          TestSignalName => "P1CMDBL(1)",
          TestDelay => tisd_P1CMDBL_P1CMDCLK(1),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBL_P1CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P1CMDBL_P1CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P1CMDBL_P1CMDCLK_negedge_posedge(1),
          HoldLow => thold_P1CMDBL_P1CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBL_P1CMDCLK_posedge(2),
          TimingData => Tmkr_P1CMDBL_P1CMDCLK_posedge(2),
          TestSignal => P1CMDBL_P1CMDCLK_dly(2),
          TestSignalName => "P1CMDBL(2)",
          TestDelay => tisd_P1CMDBL_P1CMDCLK(2),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBL_P1CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P1CMDBL_P1CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P1CMDBL_P1CMDCLK_negedge_posedge(2),
          HoldLow => thold_P1CMDBL_P1CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBL_P1CMDCLK_posedge(3),
          TimingData => Tmkr_P1CMDBL_P1CMDCLK_posedge(3),
          TestSignal => P1CMDBL_P1CMDCLK_dly(3),
          TestSignalName => "P1CMDBL(3)",
          TestDelay => tisd_P1CMDBL_P1CMDCLK(3),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBL_P1CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P1CMDBL_P1CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P1CMDBL_P1CMDCLK_negedge_posedge(3),
          HoldLow => thold_P1CMDBL_P1CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBL_P1CMDCLK_posedge(4),
          TimingData => Tmkr_P1CMDBL_P1CMDCLK_posedge(4),
          TestSignal => P1CMDBL_P1CMDCLK_dly(4),
          TestSignalName => "P1CMDBL(4)",
          TestDelay => tisd_P1CMDBL_P1CMDCLK(4),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBL_P1CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P1CMDBL_P1CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P1CMDBL_P1CMDCLK_negedge_posedge(4),
          HoldLow => thold_P1CMDBL_P1CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDBL_P1CMDCLK_posedge(5),
          TimingData => Tmkr_P1CMDBL_P1CMDCLK_posedge(5),
          TestSignal => P1CMDBL_P1CMDCLK_dly(5),
          TestSignalName => "P1CMDBL(5)",
          TestDelay => tisd_P1CMDBL_P1CMDCLK(5),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDBL_P1CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P1CMDBL_P1CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P1CMDBL_P1CMDCLK_negedge_posedge(5),
          HoldLow => thold_P1CMDBL_P1CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(0),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(0),
          TestSignal => P1CMDCA_P1CMDCLK_dly(0),
          TestSignalName => "P1CMDCA(0)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(0),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(0),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(1),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(1),
          TestSignal => P1CMDCA_P1CMDCLK_dly(1),
          TestSignalName => "P1CMDCA(1)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(1),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(1),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(10),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(10),
          TestSignal => P1CMDCA_P1CMDCLK_dly(10),
          TestSignalName => "P1CMDCA(10)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(10),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(10),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(11),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(11),
          TestSignal => P1CMDCA_P1CMDCLK_dly(11),
          TestSignalName => "P1CMDCA(11)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(11),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(11),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(2),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(2),
          TestSignal => P1CMDCA_P1CMDCLK_dly(2),
          TestSignalName => "P1CMDCA(2)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(2),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(2),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(3),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(3),
          TestSignal => P1CMDCA_P1CMDCLK_dly(3),
          TestSignalName => "P1CMDCA(3)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(3),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(3),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(4),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(4),
          TestSignal => P1CMDCA_P1CMDCLK_dly(4),
          TestSignalName => "P1CMDCA(4)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(4),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(4),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(5),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(5),
          TestSignal => P1CMDCA_P1CMDCLK_dly(5),
          TestSignalName => "P1CMDCA(5)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(5),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(5),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(6),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(6),
          TestSignal => P1CMDCA_P1CMDCLK_dly(6),
          TestSignalName => "P1CMDCA(6)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(6),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(6),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(7),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(7),
          TestSignal => P1CMDCA_P1CMDCLK_dly(7),
          TestSignalName => "P1CMDCA(7)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(7),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(7),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(8),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(8),
          TestSignal => P1CMDCA_P1CMDCLK_dly(8),
          TestSignalName => "P1CMDCA(8)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(8),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(8),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDCA_P1CMDCLK_posedge(9),
          TimingData => Tmkr_P1CMDCA_P1CMDCLK_posedge(9),
          TestSignal => P1CMDCA_P1CMDCLK_dly(9),
          TestSignalName => "P1CMDCA(9)",
          TestDelay => tisd_P1CMDCA_P1CMDCLK(9),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDCA_P1CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P1CMDCA_P1CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P1CMDCA_P1CMDCLK_negedge_posedge(9),
          HoldLow => thold_P1CMDCA_P1CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDEN_P1CMDCLK_posedge,
          TimingData => Tmkr_P1CMDEN_P1CMDCLK_posedge,
          TestSignal => P1CMDEN_P1CMDCLK_dly,
          TestSignalName => "P1CMDEN",
          TestDelay => tisd_P1CMDEN_P1CMDCLK,
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDEN_P1CMDCLK_posedge_posedge,
          HoldHigh => thold_P1CMDEN_P1CMDCLK_posedge_posedge,
          SetupLow => tsetup_P1CMDEN_P1CMDCLK_negedge_posedge,
          HoldLow => thold_P1CMDEN_P1CMDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDINSTR_P1CMDCLK_posedge(0),
          TimingData => Tmkr_P1CMDINSTR_P1CMDCLK_posedge(0),
          TestSignal => P1CMDINSTR_P1CMDCLK_dly(0),
          TestSignalName => "P1CMDINSTR(0)",
          TestDelay => tisd_P1CMDINSTR_P1CMDCLK(0),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDINSTR_P1CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P1CMDINSTR_P1CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P1CMDINSTR_P1CMDCLK_negedge_posedge(0),
          HoldLow => thold_P1CMDINSTR_P1CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDINSTR_P1CMDCLK_posedge(1),
          TimingData => Tmkr_P1CMDINSTR_P1CMDCLK_posedge(1),
          TestSignal => P1CMDINSTR_P1CMDCLK_dly(1),
          TestSignalName => "P1CMDINSTR(1)",
          TestDelay => tisd_P1CMDINSTR_P1CMDCLK(1),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDINSTR_P1CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P1CMDINSTR_P1CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P1CMDINSTR_P1CMDCLK_negedge_posedge(1),
          HoldLow => thold_P1CMDINSTR_P1CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDINSTR_P1CMDCLK_posedge(2),
          TimingData => Tmkr_P1CMDINSTR_P1CMDCLK_posedge(2),
          TestSignal => P1CMDINSTR_P1CMDCLK_dly(2),
          TestSignalName => "P1CMDINSTR(2)",
          TestDelay => tisd_P1CMDINSTR_P1CMDCLK(2),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDINSTR_P1CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P1CMDINSTR_P1CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P1CMDINSTR_P1CMDCLK_negedge_posedge(2),
          HoldLow => thold_P1CMDINSTR_P1CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(0),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(0),
          TestSignal => P1CMDRA_P1CMDCLK_dly(0),
          TestSignalName => "P1CMDRA(0)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(0),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(0),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(1),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(1),
          TestSignal => P1CMDRA_P1CMDCLK_dly(1),
          TestSignalName => "P1CMDRA(1)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(1),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(1),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(10),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(10),
          TestSignal => P1CMDRA_P1CMDCLK_dly(10),
          TestSignalName => "P1CMDRA(10)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(10),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(10),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(11),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(11),
          TestSignal => P1CMDRA_P1CMDCLK_dly(11),
          TestSignalName => "P1CMDRA(11)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(11),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(11),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(12),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(12),
          TestSignal => P1CMDRA_P1CMDCLK_dly(12),
          TestSignalName => "P1CMDRA(12)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(12),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(12),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(12),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(12),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(13),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(13),
          TestSignal => P1CMDRA_P1CMDCLK_dly(13),
          TestSignalName => "P1CMDRA(13)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(13),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(13),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(13),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(13),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(14),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(14),
          TestSignal => P1CMDRA_P1CMDCLK_dly(14),
          TestSignalName => "P1CMDRA(14)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(14),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(14),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(14),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(14),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(2),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(2),
          TestSignal => P1CMDRA_P1CMDCLK_dly(2),
          TestSignalName => "P1CMDRA(2)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(2),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(2),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(3),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(3),
          TestSignal => P1CMDRA_P1CMDCLK_dly(3),
          TestSignalName => "P1CMDRA(3)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(3),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(3),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(4),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(4),
          TestSignal => P1CMDRA_P1CMDCLK_dly(4),
          TestSignalName => "P1CMDRA(4)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(4),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(4),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(5),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(5),
          TestSignal => P1CMDRA_P1CMDCLK_dly(5),
          TestSignalName => "P1CMDRA(5)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(5),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(5),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(6),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(6),
          TestSignal => P1CMDRA_P1CMDCLK_dly(6),
          TestSignalName => "P1CMDRA(6)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(6),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(6),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(7),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(7),
          TestSignal => P1CMDRA_P1CMDCLK_dly(7),
          TestSignalName => "P1CMDRA(7)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(7),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(7),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(8),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(8),
          TestSignal => P1CMDRA_P1CMDCLK_dly(8),
          TestSignalName => "P1CMDRA(8)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(8),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(8),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1CMDRA_P1CMDCLK_posedge(9),
          TimingData => Tmkr_P1CMDRA_P1CMDCLK_posedge(9),
          TestSignal => P1CMDRA_P1CMDCLK_dly(9),
          TestSignalName => "P1CMDRA(9)",
          TestDelay => tisd_P1CMDRA_P1CMDCLK(9),
          RefSignal => P1CMDCLK_dly,
          RefSignalName => "P1CMDCLK",
          RefDelay => ticd_P1CMDCLK,
          SetupHigh => tsetup_P1CMDRA_P1CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P1CMDRA_P1CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P1CMDRA_P1CMDCLK_negedge_posedge(9),
          HoldLow => thold_P1CMDRA_P1CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1RDEN_P1RDCLK_posedge,
          TimingData => Tmkr_P1RDEN_P1RDCLK_posedge,
          TestSignal => P1RDEN_P1RDCLK_dly,
          TestSignalName => "P1RDEN",
          TestDelay => tisd_P1RDEN_P1RDCLK,
          RefSignal => P1RDCLK_dly,
          RefSignalName => "P1RDCLK",
          RefDelay => ticd_P1RDCLK,
          SetupHigh => tsetup_P1RDEN_P1RDCLK_posedge_posedge,
          HoldHigh => thold_P1RDEN_P1RDCLK_posedge_posedge,
          SetupLow => tsetup_P1RDEN_P1RDCLK_negedge_posedge,
          HoldLow => thold_P1RDEN_P1RDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1RWRMASK_P1WRCLK_posedge(0),
          TimingData => Tmkr_P1RWRMASK_P1WRCLK_posedge(0),
          TestSignal => P1RWRMASK_P1WRCLK_dly(0),
          TestSignalName => "P1RWRMASK(0)",
          TestDelay => tisd_P1RWRMASK_P1WRCLK(0),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1RWRMASK_P1WRCLK_posedge_posedge(0),
          HoldHigh => thold_P1RWRMASK_P1WRCLK_posedge_posedge(0),
          SetupLow => tsetup_P1RWRMASK_P1WRCLK_negedge_posedge(0),
          HoldLow => thold_P1RWRMASK_P1WRCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1RWRMASK_P1WRCLK_posedge(1),
          TimingData => Tmkr_P1RWRMASK_P1WRCLK_posedge(1),
          TestSignal => P1RWRMASK_P1WRCLK_dly(1),
          TestSignalName => "P1RWRMASK(1)",
          TestDelay => tisd_P1RWRMASK_P1WRCLK(1),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1RWRMASK_P1WRCLK_posedge_posedge(1),
          HoldHigh => thold_P1RWRMASK_P1WRCLK_posedge_posedge(1),
          SetupLow => tsetup_P1RWRMASK_P1WRCLK_negedge_posedge(1),
          HoldLow => thold_P1RWRMASK_P1WRCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1RWRMASK_P1WRCLK_posedge(2),
          TimingData => Tmkr_P1RWRMASK_P1WRCLK_posedge(2),
          TestSignal => P1RWRMASK_P1WRCLK_dly(2),
          TestSignalName => "P1RWRMASK(2)",
          TestDelay => tisd_P1RWRMASK_P1WRCLK(2),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1RWRMASK_P1WRCLK_posedge_posedge(2),
          HoldHigh => thold_P1RWRMASK_P1WRCLK_posedge_posedge(2),
          SetupLow => tsetup_P1RWRMASK_P1WRCLK_negedge_posedge(2),
          HoldLow => thold_P1RWRMASK_P1WRCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1RWRMASK_P1WRCLK_posedge(3),
          TimingData => Tmkr_P1RWRMASK_P1WRCLK_posedge(3),
          TestSignal => P1RWRMASK_P1WRCLK_dly(3),
          TestSignalName => "P1RWRMASK(3)",
          TestDelay => tisd_P1RWRMASK_P1WRCLK(3),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1RWRMASK_P1WRCLK_posedge_posedge(3),
          HoldHigh => thold_P1RWRMASK_P1WRCLK_posedge_posedge(3),
          SetupLow => tsetup_P1RWRMASK_P1WRCLK_negedge_posedge(3),
          HoldLow => thold_P1RWRMASK_P1WRCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(0),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(0),
          TestSignal => P1WRDATA_P1WRCLK_dly(0),
          TestSignalName => "P1WRDATA(0)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(0),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(0),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(0),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(0),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(1),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(1),
          TestSignal => P1WRDATA_P1WRCLK_dly(1),
          TestSignalName => "P1WRDATA(1)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(1),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(1),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(1),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(1),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(10),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(10),
          TestSignal => P1WRDATA_P1WRCLK_dly(10),
          TestSignalName => "P1WRDATA(10)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(10),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(10),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(10),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(10),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(11),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(11),
          TestSignal => P1WRDATA_P1WRCLK_dly(11),
          TestSignalName => "P1WRDATA(11)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(11),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(11),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(11),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(11),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(12),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(12),
          TestSignal => P1WRDATA_P1WRCLK_dly(12),
          TestSignalName => "P1WRDATA(12)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(12),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(12),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(12),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(12),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(13),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(13),
          TestSignal => P1WRDATA_P1WRCLK_dly(13),
          TestSignalName => "P1WRDATA(13)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(13),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(13),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(13),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(13),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(14),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(14),
          TestSignal => P1WRDATA_P1WRCLK_dly(14),
          TestSignalName => "P1WRDATA(14)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(14),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(14),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(14),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(14),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(15),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(15),
          TestSignal => P1WRDATA_P1WRCLK_dly(15),
          TestSignalName => "P1WRDATA(15)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(15),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(15),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(15),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(15),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(15),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(16),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(16),
          TestSignal => P1WRDATA_P1WRCLK_dly(16),
          TestSignalName => "P1WRDATA(16)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(16),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(16),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(16),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(16),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(16),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(17),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(17),
          TestSignal => P1WRDATA_P1WRCLK_dly(17),
          TestSignalName => "P1WRDATA(17)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(17),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(17),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(17),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(17),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(17),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(18),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(18),
          TestSignal => P1WRDATA_P1WRCLK_dly(18),
          TestSignalName => "P1WRDATA(18)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(18),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(18),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(18),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(18),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(18),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(19),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(19),
          TestSignal => P1WRDATA_P1WRCLK_dly(19),
          TestSignalName => "P1WRDATA(19)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(19),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(19),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(19),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(19),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(19),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(2),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(2),
          TestSignal => P1WRDATA_P1WRCLK_dly(2),
          TestSignalName => "P1WRDATA(2)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(2),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(2),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(2),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(2),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(20),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(20),
          TestSignal => P1WRDATA_P1WRCLK_dly(20),
          TestSignalName => "P1WRDATA(20)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(20),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(20),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(20),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(20),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(20),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(21),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(21),
          TestSignal => P1WRDATA_P1WRCLK_dly(21),
          TestSignalName => "P1WRDATA(21)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(21),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(21),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(21),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(21),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(21),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(22),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(22),
          TestSignal => P1WRDATA_P1WRCLK_dly(22),
          TestSignalName => "P1WRDATA(22)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(22),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(22),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(22),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(22),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(22),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(23),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(23),
          TestSignal => P1WRDATA_P1WRCLK_dly(23),
          TestSignalName => "P1WRDATA(23)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(23),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(23),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(23),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(23),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(23),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(24),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(24),
          TestSignal => P1WRDATA_P1WRCLK_dly(24),
          TestSignalName => "P1WRDATA(24)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(24),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(24),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(24),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(24),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(24),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(25),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(25),
          TestSignal => P1WRDATA_P1WRCLK_dly(25),
          TestSignalName => "P1WRDATA(25)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(25),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(25),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(25),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(25),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(25),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(26),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(26),
          TestSignal => P1WRDATA_P1WRCLK_dly(26),
          TestSignalName => "P1WRDATA(26)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(26),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(26),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(26),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(26),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(26),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(27),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(27),
          TestSignal => P1WRDATA_P1WRCLK_dly(27),
          TestSignalName => "P1WRDATA(27)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(27),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(27),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(27),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(27),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(27),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(28),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(28),
          TestSignal => P1WRDATA_P1WRCLK_dly(28),
          TestSignalName => "P1WRDATA(28)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(28),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(28),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(28),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(28),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(28),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(29),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(29),
          TestSignal => P1WRDATA_P1WRCLK_dly(29),
          TestSignalName => "P1WRDATA(29)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(29),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(29),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(29),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(29),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(29),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(3),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(3),
          TestSignal => P1WRDATA_P1WRCLK_dly(3),
          TestSignalName => "P1WRDATA(3)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(3),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(3),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(3),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(3),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(30),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(30),
          TestSignal => P1WRDATA_P1WRCLK_dly(30),
          TestSignalName => "P1WRDATA(30)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(30),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(30),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(30),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(30),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(30),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(31),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(31),
          TestSignal => P1WRDATA_P1WRCLK_dly(31),
          TestSignalName => "P1WRDATA(31)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(31),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(31),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(31),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(31),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(31),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(4),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(4),
          TestSignal => P1WRDATA_P1WRCLK_dly(4),
          TestSignalName => "P1WRDATA(4)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(4),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(4),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(4),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(4),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(5),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(5),
          TestSignal => P1WRDATA_P1WRCLK_dly(5),
          TestSignalName => "P1WRDATA(5)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(5),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(5),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(5),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(5),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(6),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(6),
          TestSignal => P1WRDATA_P1WRCLK_dly(6),
          TestSignalName => "P1WRDATA(6)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(6),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(6),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(6),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(6),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(7),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(7),
          TestSignal => P1WRDATA_P1WRCLK_dly(7),
          TestSignalName => "P1WRDATA(7)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(7),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(7),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(7),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(7),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(8),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(8),
          TestSignal => P1WRDATA_P1WRCLK_dly(8),
          TestSignalName => "P1WRDATA(8)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(8),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(8),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(8),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(8),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WRDATA_P1WRCLK_posedge(9),
          TimingData => Tmkr_P1WRDATA_P1WRCLK_posedge(9),
          TestSignal => P1WRDATA_P1WRCLK_dly(9),
          TestSignalName => "P1WRDATA(9)",
          TestDelay => tisd_P1WRDATA_P1WRCLK(9),
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WRDATA_P1WRCLK_posedge_posedge(9),
          HoldHigh => thold_P1WRDATA_P1WRCLK_posedge_posedge(9),
          SetupLow => tsetup_P1WRDATA_P1WRCLK_negedge_posedge(9),
          HoldLow => thold_P1WRDATA_P1WRCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P1WREN_P1WRCLK_posedge,
          TimingData => Tmkr_P1WREN_P1WRCLK_posedge,
          TestSignal => P1WREN_P1WRCLK_dly,
          TestSignalName => "P1WREN",
          TestDelay => tisd_P1WREN_P1WRCLK,
          RefSignal => P1WRCLK_dly,
          RefSignalName => "P1WRCLK",
          RefDelay => ticd_P1WRCLK,
          SetupHigh => tsetup_P1WREN_P1WRCLK_posedge_posedge,
          HoldHigh => thold_P1WREN_P1WRCLK_posedge_posedge,
          SetupLow => tsetup_P1WREN_P1WRCLK_negedge_posedge,
          HoldLow => thold_P1WREN_P1WRCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
         VitalSetupHoldCheck
        (
          Violation => Tviol_P2ARBEN_PLLCLK_posedge(0),
          TimingData => Tmkr_P2ARBEN_PLLCLK_posedge(0),
          TestSignal => P2ARBEN_PLLCLK_dly(0),
          TestSignalName => "P2ARBEN",
          TestDelay => tisd_P2ARBEN_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_P2ARBEN_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_P2ARBEN_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_P2ARBEN_PLLCLK_negedge_posedge(0),
          HoldLow => thold_P2ARBEN_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2ARBEN_PLLCLK_posedge(1),
          TimingData => Tmkr_P2ARBEN_PLLCLK_posedge(1),
          TestSignal => P2ARBEN_PLLCLK_dly(1),
          TestSignalName => "P2ARBEN",
          TestDelay => tisd_P2ARBEN_PLLCLK(1),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_P2ARBEN_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_P2ARBEN_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_P2ARBEN_PLLCLK_negedge_posedge(1),
          HoldLow => thold_P2ARBEN_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBA_P2CMDCLK_posedge(0),
          TimingData => Tmkr_P2CMDBA_P2CMDCLK_posedge(0),
          TestSignal => P2CMDBA_P2CMDCLK_dly(0),
          TestSignalName => "P2CMDBA(0)",
          TestDelay => tisd_P2CMDBA_P2CMDCLK(0),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBA_P2CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P2CMDBA_P2CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P2CMDBA_P2CMDCLK_negedge_posedge(0),
          HoldLow => thold_P2CMDBA_P2CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBA_P2CMDCLK_posedge(1),
          TimingData => Tmkr_P2CMDBA_P2CMDCLK_posedge(1),
          TestSignal => P2CMDBA_P2CMDCLK_dly(1),
          TestSignalName => "P2CMDBA(1)",
          TestDelay => tisd_P2CMDBA_P2CMDCLK(1),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBA_P2CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P2CMDBA_P2CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P2CMDBA_P2CMDCLK_negedge_posedge(1),
          HoldLow => thold_P2CMDBA_P2CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBA_P2CMDCLK_posedge(2),
          TimingData => Tmkr_P2CMDBA_P2CMDCLK_posedge(2),
          TestSignal => P2CMDBA_P2CMDCLK_dly(2),
          TestSignalName => "P2CMDBA(2)",
          TestDelay => tisd_P2CMDBA_P2CMDCLK(2),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBA_P2CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P2CMDBA_P2CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P2CMDBA_P2CMDCLK_negedge_posedge(2),
          HoldLow => thold_P2CMDBA_P2CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBL_P2CMDCLK_posedge(0),
          TimingData => Tmkr_P2CMDBL_P2CMDCLK_posedge(0),
          TestSignal => P2CMDBL_P2CMDCLK_dly(0),
          TestSignalName => "P2CMDBL(0)",
          TestDelay => tisd_P2CMDBL_P2CMDCLK(0),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBL_P2CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P2CMDBL_P2CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P2CMDBL_P2CMDCLK_negedge_posedge(0),
          HoldLow => thold_P2CMDBL_P2CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBL_P2CMDCLK_posedge(1),
          TimingData => Tmkr_P2CMDBL_P2CMDCLK_posedge(1),
          TestSignal => P2CMDBL_P2CMDCLK_dly(1),
          TestSignalName => "P2CMDBL(1)",
          TestDelay => tisd_P2CMDBL_P2CMDCLK(1),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBL_P2CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P2CMDBL_P2CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P2CMDBL_P2CMDCLK_negedge_posedge(1),
          HoldLow => thold_P2CMDBL_P2CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBL_P2CMDCLK_posedge(2),
          TimingData => Tmkr_P2CMDBL_P2CMDCLK_posedge(2),
          TestSignal => P2CMDBL_P2CMDCLK_dly(2),
          TestSignalName => "P2CMDBL(2)",
          TestDelay => tisd_P2CMDBL_P2CMDCLK(2),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBL_P2CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P2CMDBL_P2CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P2CMDBL_P2CMDCLK_negedge_posedge(2),
          HoldLow => thold_P2CMDBL_P2CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBL_P2CMDCLK_posedge(3),
          TimingData => Tmkr_P2CMDBL_P2CMDCLK_posedge(3),
          TestSignal => P2CMDBL_P2CMDCLK_dly(3),
          TestSignalName => "P2CMDBL(3)",
          TestDelay => tisd_P2CMDBL_P2CMDCLK(3),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBL_P2CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P2CMDBL_P2CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P2CMDBL_P2CMDCLK_negedge_posedge(3),
          HoldLow => thold_P2CMDBL_P2CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBL_P2CMDCLK_posedge(4),
          TimingData => Tmkr_P2CMDBL_P2CMDCLK_posedge(4),
          TestSignal => P2CMDBL_P2CMDCLK_dly(4),
          TestSignalName => "P2CMDBL(4)",
          TestDelay => tisd_P2CMDBL_P2CMDCLK(4),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBL_P2CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P2CMDBL_P2CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P2CMDBL_P2CMDCLK_negedge_posedge(4),
          HoldLow => thold_P2CMDBL_P2CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDBL_P2CMDCLK_posedge(5),
          TimingData => Tmkr_P2CMDBL_P2CMDCLK_posedge(5),
          TestSignal => P2CMDBL_P2CMDCLK_dly(5),
          TestSignalName => "P2CMDBL(5)",
          TestDelay => tisd_P2CMDBL_P2CMDCLK(5),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDBL_P2CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P2CMDBL_P2CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P2CMDBL_P2CMDCLK_negedge_posedge(5),
          HoldLow => thold_P2CMDBL_P2CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(0),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(0),
          TestSignal => P2CMDCA_P2CMDCLK_dly(0),
          TestSignalName => "P2CMDCA(0)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(0),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(0),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(1),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(1),
          TestSignal => P2CMDCA_P2CMDCLK_dly(1),
          TestSignalName => "P2CMDCA(1)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(1),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(1),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(10),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(10),
          TestSignal => P2CMDCA_P2CMDCLK_dly(10),
          TestSignalName => "P2CMDCA(10)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(10),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(10),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(11),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(11),
          TestSignal => P2CMDCA_P2CMDCLK_dly(11),
          TestSignalName => "P2CMDCA(11)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(11),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(11),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(2),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(2),
          TestSignal => P2CMDCA_P2CMDCLK_dly(2),
          TestSignalName => "P2CMDCA(2)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(2),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(2),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(3),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(3),
          TestSignal => P2CMDCA_P2CMDCLK_dly(3),
          TestSignalName => "P2CMDCA(3)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(3),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(3),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(4),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(4),
          TestSignal => P2CMDCA_P2CMDCLK_dly(4),
          TestSignalName => "P2CMDCA(4)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(4),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(4),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(5),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(5),
          TestSignal => P2CMDCA_P2CMDCLK_dly(5),
          TestSignalName => "P2CMDCA(5)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(5),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(5),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(6),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(6),
          TestSignal => P2CMDCA_P2CMDCLK_dly(6),
          TestSignalName => "P2CMDCA(6)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(6),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(6),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(7),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(7),
          TestSignal => P2CMDCA_P2CMDCLK_dly(7),
          TestSignalName => "P2CMDCA(7)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(7),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(7),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(8),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(8),
          TestSignal => P2CMDCA_P2CMDCLK_dly(8),
          TestSignalName => "P2CMDCA(8)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(8),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(8),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDCA_P2CMDCLK_posedge(9),
          TimingData => Tmkr_P2CMDCA_P2CMDCLK_posedge(9),
          TestSignal => P2CMDCA_P2CMDCLK_dly(9),
          TestSignalName => "P2CMDCA(9)",
          TestDelay => tisd_P2CMDCA_P2CMDCLK(9),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDCA_P2CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P2CMDCA_P2CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P2CMDCA_P2CMDCLK_negedge_posedge(9),
          HoldLow => thold_P2CMDCA_P2CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDEN_P2CMDCLK_posedge,
          TimingData => Tmkr_P2CMDEN_P2CMDCLK_posedge,
          TestSignal => P2CMDEN_P2CMDCLK_dly,
          TestSignalName => "P2CMDEN",
          TestDelay => tisd_P2CMDEN_P2CMDCLK,
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDEN_P2CMDCLK_posedge_posedge,
          HoldHigh => thold_P2CMDEN_P2CMDCLK_posedge_posedge,
          SetupLow => tsetup_P2CMDEN_P2CMDCLK_negedge_posedge,
          HoldLow => thold_P2CMDEN_P2CMDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDINSTR_P2CMDCLK_posedge(0),
          TimingData => Tmkr_P2CMDINSTR_P2CMDCLK_posedge(0),
          TestSignal => P2CMDINSTR_P2CMDCLK_dly(0),
          TestSignalName => "P2CMDINSTR(0)",
          TestDelay => tisd_P2CMDINSTR_P2CMDCLK(0),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDINSTR_P2CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P2CMDINSTR_P2CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P2CMDINSTR_P2CMDCLK_negedge_posedge(0),
          HoldLow => thold_P2CMDINSTR_P2CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDINSTR_P2CMDCLK_posedge(1),
          TimingData => Tmkr_P2CMDINSTR_P2CMDCLK_posedge(1),
          TestSignal => P2CMDINSTR_P2CMDCLK_dly(1),
          TestSignalName => "P2CMDINSTR(1)",
          TestDelay => tisd_P2CMDINSTR_P2CMDCLK(1),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDINSTR_P2CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P2CMDINSTR_P2CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P2CMDINSTR_P2CMDCLK_negedge_posedge(1),
          HoldLow => thold_P2CMDINSTR_P2CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDINSTR_P2CMDCLK_posedge(2),
          TimingData => Tmkr_P2CMDINSTR_P2CMDCLK_posedge(2),
          TestSignal => P2CMDINSTR_P2CMDCLK_dly(2),
          TestSignalName => "P2CMDINSTR(2)",
          TestDelay => tisd_P2CMDINSTR_P2CMDCLK(2),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDINSTR_P2CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P2CMDINSTR_P2CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P2CMDINSTR_P2CMDCLK_negedge_posedge(2),
          HoldLow => thold_P2CMDINSTR_P2CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(0),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(0),
          TestSignal => P2CMDRA_P2CMDCLK_dly(0),
          TestSignalName => "P2CMDRA(0)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(0),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(0),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(1),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(1),
          TestSignal => P2CMDRA_P2CMDCLK_dly(1),
          TestSignalName => "P2CMDRA(1)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(1),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(1),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(10),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(10),
          TestSignal => P2CMDRA_P2CMDCLK_dly(10),
          TestSignalName => "P2CMDRA(10)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(10),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(10),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(11),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(11),
          TestSignal => P2CMDRA_P2CMDCLK_dly(11),
          TestSignalName => "P2CMDRA(11)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(11),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(11),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(12),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(12),
          TestSignal => P2CMDRA_P2CMDCLK_dly(12),
          TestSignalName => "P2CMDRA(12)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(12),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(12),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(12),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(12),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(13),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(13),
          TestSignal => P2CMDRA_P2CMDCLK_dly(13),
          TestSignalName => "P2CMDRA(13)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(13),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(13),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(13),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(13),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(14),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(14),
          TestSignal => P2CMDRA_P2CMDCLK_dly(14),
          TestSignalName => "P2CMDRA(14)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(14),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(14),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(14),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(14),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(2),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(2),
          TestSignal => P2CMDRA_P2CMDCLK_dly(2),
          TestSignalName => "P2CMDRA(2)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(2),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(2),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(3),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(3),
          TestSignal => P2CMDRA_P2CMDCLK_dly(3),
          TestSignalName => "P2CMDRA(3)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(3),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(3),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(4),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(4),
          TestSignal => P2CMDRA_P2CMDCLK_dly(4),
          TestSignalName => "P2CMDRA(4)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(4),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(4),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(5),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(5),
          TestSignal => P2CMDRA_P2CMDCLK_dly(5),
          TestSignalName => "P2CMDRA(5)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(5),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(5),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(6),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(6),
          TestSignal => P2CMDRA_P2CMDCLK_dly(6),
          TestSignalName => "P2CMDRA(6)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(6),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(6),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(7),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(7),
          TestSignal => P2CMDRA_P2CMDCLK_dly(7),
          TestSignalName => "P2CMDRA(7)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(7),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(7),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(8),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(8),
          TestSignal => P2CMDRA_P2CMDCLK_dly(8),
          TestSignalName => "P2CMDRA(8)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(8),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(8),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2CMDRA_P2CMDCLK_posedge(9),
          TimingData => Tmkr_P2CMDRA_P2CMDCLK_posedge(9),
          TestSignal => P2CMDRA_P2CMDCLK_dly(9),
          TestSignalName => "P2CMDRA(9)",
          TestDelay => tisd_P2CMDRA_P2CMDCLK(9),
          RefSignal => P2CMDCLK_dly,
          RefSignalName => "P2CMDCLK",
          RefDelay => ticd_P2CMDCLK,
          SetupHigh => tsetup_P2CMDRA_P2CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P2CMDRA_P2CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P2CMDRA_P2CMDCLK_negedge_posedge(9),
          HoldLow => thold_P2CMDRA_P2CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2EN_P2CLK_posedge,
          TimingData => Tmkr_P2EN_P2CLK_posedge,
          TestSignal => P2EN_P2CLK_dly,
          TestSignalName => "P2EN",
          TestDelay => tisd_P2EN_P2CLK,
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2EN_P2CLK_posedge_posedge,
          HoldHigh => thold_P2EN_P2CLK_posedge_posedge,
          SetupLow => tsetup_P2EN_P2CLK_negedge_posedge,
          HoldLow => thold_P2EN_P2CLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(0),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(0),
          TestSignal => P2WRDATA_P2CLK_dly(0),
          TestSignalName => "P2WRDATA(0)",
          TestDelay => tisd_P2WRDATA_P2CLK(0),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(0),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(0),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(0),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(1),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(1),
          TestSignal => P2WRDATA_P2CLK_dly(1),
          TestSignalName => "P2WRDATA(1)",
          TestDelay => tisd_P2WRDATA_P2CLK(1),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(1),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(1),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(1),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(10),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(10),
          TestSignal => P2WRDATA_P2CLK_dly(10),
          TestSignalName => "P2WRDATA(10)",
          TestDelay => tisd_P2WRDATA_P2CLK(10),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(10),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(10),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(10),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(11),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(11),
          TestSignal => P2WRDATA_P2CLK_dly(11),
          TestSignalName => "P2WRDATA(11)",
          TestDelay => tisd_P2WRDATA_P2CLK(11),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(11),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(11),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(11),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(12),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(12),
          TestSignal => P2WRDATA_P2CLK_dly(12),
          TestSignalName => "P2WRDATA(12)",
          TestDelay => tisd_P2WRDATA_P2CLK(12),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(12),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(12),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(12),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(13),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(13),
          TestSignal => P2WRDATA_P2CLK_dly(13),
          TestSignalName => "P2WRDATA(13)",
          TestDelay => tisd_P2WRDATA_P2CLK(13),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(13),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(13),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(13),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(14),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(14),
          TestSignal => P2WRDATA_P2CLK_dly(14),
          TestSignalName => "P2WRDATA(14)",
          TestDelay => tisd_P2WRDATA_P2CLK(14),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(14),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(14),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(14),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(15),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(15),
          TestSignal => P2WRDATA_P2CLK_dly(15),
          TestSignalName => "P2WRDATA(15)",
          TestDelay => tisd_P2WRDATA_P2CLK(15),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(15),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(15),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(15),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(15),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(16),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(16),
          TestSignal => P2WRDATA_P2CLK_dly(16),
          TestSignalName => "P2WRDATA(16)",
          TestDelay => tisd_P2WRDATA_P2CLK(16),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(16),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(16),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(16),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(16),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(17),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(17),
          TestSignal => P2WRDATA_P2CLK_dly(17),
          TestSignalName => "P2WRDATA(17)",
          TestDelay => tisd_P2WRDATA_P2CLK(17),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(17),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(17),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(17),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(17),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(18),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(18),
          TestSignal => P2WRDATA_P2CLK_dly(18),
          TestSignalName => "P2WRDATA(18)",
          TestDelay => tisd_P2WRDATA_P2CLK(18),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(18),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(18),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(18),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(18),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(19),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(19),
          TestSignal => P2WRDATA_P2CLK_dly(19),
          TestSignalName => "P2WRDATA(19)",
          TestDelay => tisd_P2WRDATA_P2CLK(19),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(19),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(19),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(19),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(19),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(2),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(2),
          TestSignal => P2WRDATA_P2CLK_dly(2),
          TestSignalName => "P2WRDATA(2)",
          TestDelay => tisd_P2WRDATA_P2CLK(2),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(2),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(2),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(2),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(20),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(20),
          TestSignal => P2WRDATA_P2CLK_dly(20),
          TestSignalName => "P2WRDATA(20)",
          TestDelay => tisd_P2WRDATA_P2CLK(20),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(20),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(20),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(20),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(20),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(21),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(21),
          TestSignal => P2WRDATA_P2CLK_dly(21),
          TestSignalName => "P2WRDATA(21)",
          TestDelay => tisd_P2WRDATA_P2CLK(21),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(21),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(21),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(21),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(21),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(22),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(22),
          TestSignal => P2WRDATA_P2CLK_dly(22),
          TestSignalName => "P2WRDATA(22)",
          TestDelay => tisd_P2WRDATA_P2CLK(22),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(22),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(22),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(22),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(22),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(23),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(23),
          TestSignal => P2WRDATA_P2CLK_dly(23),
          TestSignalName => "P2WRDATA(23)",
          TestDelay => tisd_P2WRDATA_P2CLK(23),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(23),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(23),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(23),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(23),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(24),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(24),
          TestSignal => P2WRDATA_P2CLK_dly(24),
          TestSignalName => "P2WRDATA(24)",
          TestDelay => tisd_P2WRDATA_P2CLK(24),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(24),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(24),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(24),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(24),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(25),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(25),
          TestSignal => P2WRDATA_P2CLK_dly(25),
          TestSignalName => "P2WRDATA(25)",
          TestDelay => tisd_P2WRDATA_P2CLK(25),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(25),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(25),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(25),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(25),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(26),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(26),
          TestSignal => P2WRDATA_P2CLK_dly(26),
          TestSignalName => "P2WRDATA(26)",
          TestDelay => tisd_P2WRDATA_P2CLK(26),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(26),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(26),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(26),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(26),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(27),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(27),
          TestSignal => P2WRDATA_P2CLK_dly(27),
          TestSignalName => "P2WRDATA(27)",
          TestDelay => tisd_P2WRDATA_P2CLK(27),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(27),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(27),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(27),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(27),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(28),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(28),
          TestSignal => P2WRDATA_P2CLK_dly(28),
          TestSignalName => "P2WRDATA(28)",
          TestDelay => tisd_P2WRDATA_P2CLK(28),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(28),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(28),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(28),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(28),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(29),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(29),
          TestSignal => P2WRDATA_P2CLK_dly(29),
          TestSignalName => "P2WRDATA(29)",
          TestDelay => tisd_P2WRDATA_P2CLK(29),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(29),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(29),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(29),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(29),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(3),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(3),
          TestSignal => P2WRDATA_P2CLK_dly(3),
          TestSignalName => "P2WRDATA(3)",
          TestDelay => tisd_P2WRDATA_P2CLK(3),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(3),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(3),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(3),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(30),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(30),
          TestSignal => P2WRDATA_P2CLK_dly(30),
          TestSignalName => "P2WRDATA(30)",
          TestDelay => tisd_P2WRDATA_P2CLK(30),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(30),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(30),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(30),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(30),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(31),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(31),
          TestSignal => P2WRDATA_P2CLK_dly(31),
          TestSignalName => "P2WRDATA(31)",
          TestDelay => tisd_P2WRDATA_P2CLK(31),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(31),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(31),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(31),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(31),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(4),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(4),
          TestSignal => P2WRDATA_P2CLK_dly(4),
          TestSignalName => "P2WRDATA(4)",
          TestDelay => tisd_P2WRDATA_P2CLK(4),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(4),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(4),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(4),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(5),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(5),
          TestSignal => P2WRDATA_P2CLK_dly(5),
          TestSignalName => "P2WRDATA(5)",
          TestDelay => tisd_P2WRDATA_P2CLK(5),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(5),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(5),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(5),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(6),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(6),
          TestSignal => P2WRDATA_P2CLK_dly(6),
          TestSignalName => "P2WRDATA(6)",
          TestDelay => tisd_P2WRDATA_P2CLK(6),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(6),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(6),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(6),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(7),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(7),
          TestSignal => P2WRDATA_P2CLK_dly(7),
          TestSignalName => "P2WRDATA(7)",
          TestDelay => tisd_P2WRDATA_P2CLK(7),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(7),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(7),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(7),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(8),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(8),
          TestSignal => P2WRDATA_P2CLK_dly(8),
          TestSignalName => "P2WRDATA(8)",
          TestDelay => tisd_P2WRDATA_P2CLK(8),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(8),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(8),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(8),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRDATA_P2CLK_posedge(9),
          TimingData => Tmkr_P2WRDATA_P2CLK_posedge(9),
          TestSignal => P2WRDATA_P2CLK_dly(9),
          TestSignalName => "P2WRDATA(9)",
          TestDelay => tisd_P2WRDATA_P2CLK(9),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRDATA_P2CLK_posedge_posedge(9),
          HoldHigh => thold_P2WRDATA_P2CLK_posedge_posedge(9),
          SetupLow => tsetup_P2WRDATA_P2CLK_negedge_posedge(9),
          HoldLow => thold_P2WRDATA_P2CLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRMASK_P2CLK_posedge(0),
          TimingData => Tmkr_P2WRMASK_P2CLK_posedge(0),
          TestSignal => P2WRMASK_P2CLK_dly(0),
          TestSignalName => "P2WRMASK(0)",
          TestDelay => tisd_P2WRMASK_P2CLK(0),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRMASK_P2CLK_posedge_posedge(0),
          HoldHigh => thold_P2WRMASK_P2CLK_posedge_posedge(0),
          SetupLow => tsetup_P2WRMASK_P2CLK_negedge_posedge(0),
          HoldLow => thold_P2WRMASK_P2CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRMASK_P2CLK_posedge(1),
          TimingData => Tmkr_P2WRMASK_P2CLK_posedge(1),
          TestSignal => P2WRMASK_P2CLK_dly(1),
          TestSignalName => "P2WRMASK(1)",
          TestDelay => tisd_P2WRMASK_P2CLK(1),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRMASK_P2CLK_posedge_posedge(1),
          HoldHigh => thold_P2WRMASK_P2CLK_posedge_posedge(1),
          SetupLow => tsetup_P2WRMASK_P2CLK_negedge_posedge(1),
          HoldLow => thold_P2WRMASK_P2CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRMASK_P2CLK_posedge(2),
          TimingData => Tmkr_P2WRMASK_P2CLK_posedge(2),
          TestSignal => P2WRMASK_P2CLK_dly(2),
          TestSignalName => "P2WRMASK(2)",
          TestDelay => tisd_P2WRMASK_P2CLK(2),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRMASK_P2CLK_posedge_posedge(2),
          HoldHigh => thold_P2WRMASK_P2CLK_posedge_posedge(2),
          SetupLow => tsetup_P2WRMASK_P2CLK_negedge_posedge(2),
          HoldLow => thold_P2WRMASK_P2CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P2WRMASK_P2CLK_posedge(3),
          TimingData => Tmkr_P2WRMASK_P2CLK_posedge(3),
          TestSignal => P2WRMASK_P2CLK_dly(3),
          TestSignalName => "P2WRMASK(3)",
          TestDelay => tisd_P2WRMASK_P2CLK(3),
          RefSignal => P2CLK_dly,
          RefSignalName => "P2CLK",
          RefDelay => ticd_P2CLK,
          SetupHigh => tsetup_P2WRMASK_P2CLK_posedge_posedge(3),
          HoldHigh => thold_P2WRMASK_P2CLK_posedge_posedge(3),
          SetupLow => tsetup_P2WRMASK_P2CLK_negedge_posedge(3),
          HoldLow => thold_P2WRMASK_P2CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3ARBEN_PLLCLK_posedge(0),
          TimingData => Tmkr_P3ARBEN_PLLCLK_posedge(0),
          TestSignal => P3ARBEN_PLLCLK_dly(0),
          TestSignalName => "P3ARBEN",
          TestDelay => tisd_P3ARBEN_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_P3ARBEN_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_P3ARBEN_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_P3ARBEN_PLLCLK_negedge_posedge(0),
          HoldLow => thold_P3ARBEN_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3ARBEN_PLLCLK_posedge(1),
          TimingData => Tmkr_P3ARBEN_PLLCLK_posedge(1),
          TestSignal => P3ARBEN_PLLCLK_dly(1),
          TestSignalName => "P3ARBEN",
          TestDelay => tisd_P3ARBEN_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_P3ARBEN_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_P3ARBEN_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_P3ARBEN_PLLCLK_negedge_posedge(1),
          HoldLow => thold_P3ARBEN_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBA_P3CMDCLK_posedge(0),
          TimingData => Tmkr_P3CMDBA_P3CMDCLK_posedge(0),
          TestSignal => P3CMDBA_P3CMDCLK_dly(0),
          TestSignalName => "P3CMDBA(0)",
          TestDelay => tisd_P3CMDBA_P3CMDCLK(0),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBA_P3CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P3CMDBA_P3CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P3CMDBA_P3CMDCLK_negedge_posedge(0),
          HoldLow => thold_P3CMDBA_P3CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBA_P3CMDCLK_posedge(1),
          TimingData => Tmkr_P3CMDBA_P3CMDCLK_posedge(1),
          TestSignal => P3CMDBA_P3CMDCLK_dly(1),
          TestSignalName => "P3CMDBA(1)",
          TestDelay => tisd_P3CMDBA_P3CMDCLK(1),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBA_P3CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P3CMDBA_P3CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P3CMDBA_P3CMDCLK_negedge_posedge(1),
          HoldLow => thold_P3CMDBA_P3CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBA_P3CMDCLK_posedge(2),
          TimingData => Tmkr_P3CMDBA_P3CMDCLK_posedge(2),
          TestSignal => P3CMDBA_P3CMDCLK_dly(2),
          TestSignalName => "P3CMDBA(2)",
          TestDelay => tisd_P3CMDBA_P3CMDCLK(2),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBA_P3CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P3CMDBA_P3CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P3CMDBA_P3CMDCLK_negedge_posedge(2),
          HoldLow => thold_P3CMDBA_P3CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBL_P3CMDCLK_posedge(0),
          TimingData => Tmkr_P3CMDBL_P3CMDCLK_posedge(0),
          TestSignal => P3CMDBL_P3CMDCLK_dly(0),
          TestSignalName => "P3CMDBL(0)",
          TestDelay => tisd_P3CMDBL_P3CMDCLK(0),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBL_P3CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P3CMDBL_P3CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P3CMDBL_P3CMDCLK_negedge_posedge(0),
          HoldLow => thold_P3CMDBL_P3CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBL_P3CMDCLK_posedge(1),
          TimingData => Tmkr_P3CMDBL_P3CMDCLK_posedge(1),
          TestSignal => P3CMDBL_P3CMDCLK_dly(1),
          TestSignalName => "P3CMDBL(1)",
          TestDelay => tisd_P3CMDBL_P3CMDCLK(1),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBL_P3CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P3CMDBL_P3CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P3CMDBL_P3CMDCLK_negedge_posedge(1),
          HoldLow => thold_P3CMDBL_P3CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBL_P3CMDCLK_posedge(2),
          TimingData => Tmkr_P3CMDBL_P3CMDCLK_posedge(2),
          TestSignal => P3CMDBL_P3CMDCLK_dly(2),
          TestSignalName => "P3CMDBL(2)",
          TestDelay => tisd_P3CMDBL_P3CMDCLK(2),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBL_P3CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P3CMDBL_P3CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P3CMDBL_P3CMDCLK_negedge_posedge(2),
          HoldLow => thold_P3CMDBL_P3CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBL_P3CMDCLK_posedge(3),
          TimingData => Tmkr_P3CMDBL_P3CMDCLK_posedge(3),
          TestSignal => P3CMDBL_P3CMDCLK_dly(3),
          TestSignalName => "P3CMDBL(3)",
          TestDelay => tisd_P3CMDBL_P3CMDCLK(3),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBL_P3CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P3CMDBL_P3CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P3CMDBL_P3CMDCLK_negedge_posedge(3),
          HoldLow => thold_P3CMDBL_P3CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBL_P3CMDCLK_posedge(4),
          TimingData => Tmkr_P3CMDBL_P3CMDCLK_posedge(4),
          TestSignal => P3CMDBL_P3CMDCLK_dly(4),
          TestSignalName => "P3CMDBL(4)",
          TestDelay => tisd_P3CMDBL_P3CMDCLK(4),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBL_P3CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P3CMDBL_P3CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P3CMDBL_P3CMDCLK_negedge_posedge(4),
          HoldLow => thold_P3CMDBL_P3CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDBL_P3CMDCLK_posedge(5),
          TimingData => Tmkr_P3CMDBL_P3CMDCLK_posedge(5),
          TestSignal => P3CMDBL_P3CMDCLK_dly(5),
          TestSignalName => "P3CMDBL(5)",
          TestDelay => tisd_P3CMDBL_P3CMDCLK(5),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDBL_P3CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P3CMDBL_P3CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P3CMDBL_P3CMDCLK_negedge_posedge(5),
          HoldLow => thold_P3CMDBL_P3CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(0),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(0),
          TestSignal => P3CMDCA_P3CMDCLK_dly(0),
          TestSignalName => "P3CMDCA(0)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(0),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(0),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(1),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(1),
          TestSignal => P3CMDCA_P3CMDCLK_dly(1),
          TestSignalName => "P3CMDCA(1)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(1),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(1),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(10),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(10),
          TestSignal => P3CMDCA_P3CMDCLK_dly(10),
          TestSignalName => "P3CMDCA(10)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(10),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(10),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(11),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(11),
          TestSignal => P3CMDCA_P3CMDCLK_dly(11),
          TestSignalName => "P3CMDCA(11)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(11),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(11),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(2),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(2),
          TestSignal => P3CMDCA_P3CMDCLK_dly(2),
          TestSignalName => "P3CMDCA(2)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(2),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(2),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(3),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(3),
          TestSignal => P3CMDCA_P3CMDCLK_dly(3),
          TestSignalName => "P3CMDCA(3)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(3),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(3),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(4),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(4),
          TestSignal => P3CMDCA_P3CMDCLK_dly(4),
          TestSignalName => "P3CMDCA(4)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(4),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(4),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(5),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(5),
          TestSignal => P3CMDCA_P3CMDCLK_dly(5),
          TestSignalName => "P3CMDCA(5)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(5),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(5),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(6),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(6),
          TestSignal => P3CMDCA_P3CMDCLK_dly(6),
          TestSignalName => "P3CMDCA(6)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(6),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(6),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(7),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(7),
          TestSignal => P3CMDCA_P3CMDCLK_dly(7),
          TestSignalName => "P3CMDCA(7)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(7),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(7),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(8),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(8),
          TestSignal => P3CMDCA_P3CMDCLK_dly(8),
          TestSignalName => "P3CMDCA(8)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(8),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(8),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDCA_P3CMDCLK_posedge(9),
          TimingData => Tmkr_P3CMDCA_P3CMDCLK_posedge(9),
          TestSignal => P3CMDCA_P3CMDCLK_dly(9),
          TestSignalName => "P3CMDCA(9)",
          TestDelay => tisd_P3CMDCA_P3CMDCLK(9),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDCA_P3CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P3CMDCA_P3CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P3CMDCA_P3CMDCLK_negedge_posedge(9),
          HoldLow => thold_P3CMDCA_P3CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDEN_P3CMDCLK_posedge,
          TimingData => Tmkr_P3CMDEN_P3CMDCLK_posedge,
          TestSignal => P3CMDEN_P3CMDCLK_dly,
          TestSignalName => "P3CMDEN",
          TestDelay => tisd_P3CMDEN_P3CMDCLK,
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDEN_P3CMDCLK_posedge_posedge,
          HoldHigh => thold_P3CMDEN_P3CMDCLK_posedge_posedge,
          SetupLow => tsetup_P3CMDEN_P3CMDCLK_negedge_posedge,
          HoldLow => thold_P3CMDEN_P3CMDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDINSTR_P3CMDCLK_posedge(0),
          TimingData => Tmkr_P3CMDINSTR_P3CMDCLK_posedge(0),
          TestSignal => P3CMDINSTR_P3CMDCLK_dly(0),
          TestSignalName => "P3CMDINSTR(0)",
          TestDelay => tisd_P3CMDINSTR_P3CMDCLK(0),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDINSTR_P3CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P3CMDINSTR_P3CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P3CMDINSTR_P3CMDCLK_negedge_posedge(0),
          HoldLow => thold_P3CMDINSTR_P3CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDINSTR_P3CMDCLK_posedge(1),
          TimingData => Tmkr_P3CMDINSTR_P3CMDCLK_posedge(1),
          TestSignal => P3CMDINSTR_P3CMDCLK_dly(1),
          TestSignalName => "P3CMDINSTR(1)",
          TestDelay => tisd_P3CMDINSTR_P3CMDCLK(1),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDINSTR_P3CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P3CMDINSTR_P3CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P3CMDINSTR_P3CMDCLK_negedge_posedge(1),
          HoldLow => thold_P3CMDINSTR_P3CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDINSTR_P3CMDCLK_posedge(2),
          TimingData => Tmkr_P3CMDINSTR_P3CMDCLK_posedge(2),
          TestSignal => P3CMDINSTR_P3CMDCLK_dly(2),
          TestSignalName => "P3CMDINSTR(2)",
          TestDelay => tisd_P3CMDINSTR_P3CMDCLK(2),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDINSTR_P3CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P3CMDINSTR_P3CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P3CMDINSTR_P3CMDCLK_negedge_posedge(2),
          HoldLow => thold_P3CMDINSTR_P3CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(0),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(0),
          TestSignal => P3CMDRA_P3CMDCLK_dly(0),
          TestSignalName => "P3CMDRA(0)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(0),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(0),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(1),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(1),
          TestSignal => P3CMDRA_P3CMDCLK_dly(1),
          TestSignalName => "P3CMDRA(1)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(1),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(1),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(10),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(10),
          TestSignal => P3CMDRA_P3CMDCLK_dly(10),
          TestSignalName => "P3CMDRA(10)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(10),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(10),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(11),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(11),
          TestSignal => P3CMDRA_P3CMDCLK_dly(11),
          TestSignalName => "P3CMDRA(11)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(11),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(11),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(12),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(12),
          TestSignal => P3CMDRA_P3CMDCLK_dly(12),
          TestSignalName => "P3CMDRA(12)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(12),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(12),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(12),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(12),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(13),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(13),
          TestSignal => P3CMDRA_P3CMDCLK_dly(13),
          TestSignalName => "P3CMDRA(13)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(13),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(13),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(13),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(13),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(14),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(14),
          TestSignal => P3CMDRA_P3CMDCLK_dly(14),
          TestSignalName => "P3CMDRA(14)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(14),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(14),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(14),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(14),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(2),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(2),
          TestSignal => P3CMDRA_P3CMDCLK_dly(2),
          TestSignalName => "P3CMDRA(2)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(2),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(2),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(3),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(3),
          TestSignal => P3CMDRA_P3CMDCLK_dly(3),
          TestSignalName => "P3CMDRA(3)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(3),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(3),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(4),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(4),
          TestSignal => P3CMDRA_P3CMDCLK_dly(4),
          TestSignalName => "P3CMDRA(4)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(4),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(4),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(5),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(5),
          TestSignal => P3CMDRA_P3CMDCLK_dly(5),
          TestSignalName => "P3CMDRA(5)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(5),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(5),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(6),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(6),
          TestSignal => P3CMDRA_P3CMDCLK_dly(6),
          TestSignalName => "P3CMDRA(6)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(6),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(6),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(7),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(7),
          TestSignal => P3CMDRA_P3CMDCLK_dly(7),
          TestSignalName => "P3CMDRA(7)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(7),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(7),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(8),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(8),
          TestSignal => P3CMDRA_P3CMDCLK_dly(8),
          TestSignalName => "P3CMDRA(8)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(8),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(8),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3CMDRA_P3CMDCLK_posedge(9),
          TimingData => Tmkr_P3CMDRA_P3CMDCLK_posedge(9),
          TestSignal => P3CMDRA_P3CMDCLK_dly(9),
          TestSignalName => "P3CMDRA(9)",
          TestDelay => tisd_P3CMDRA_P3CMDCLK(9),
          RefSignal => P3CMDCLK_dly,
          RefSignalName => "P3CMDCLK",
          RefDelay => ticd_P3CMDCLK,
          SetupHigh => tsetup_P3CMDRA_P3CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P3CMDRA_P3CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P3CMDRA_P3CMDCLK_negedge_posedge(9),
          HoldLow => thold_P3CMDRA_P3CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3EN_P3CLK_posedge,
          TimingData => Tmkr_P3EN_P3CLK_posedge,
          TestSignal => P3EN_P3CLK_dly,
          TestSignalName => "P3EN",
          TestDelay => tisd_P3EN_P3CLK,
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3EN_P3CLK_posedge_posedge,
          HoldHigh => thold_P3EN_P3CLK_posedge_posedge,
          SetupLow => tsetup_P3EN_P3CLK_negedge_posedge,
          HoldLow => thold_P3EN_P3CLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(0),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(0),
          TestSignal => P3WRDATA_P3CLK_dly(0),
          TestSignalName => "P3WRDATA(0)",
          TestDelay => tisd_P3WRDATA_P3CLK(0),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(0),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(0),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(0),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(1),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(1),
          TestSignal => P3WRDATA_P3CLK_dly(1),
          TestSignalName => "P3WRDATA(1)",
          TestDelay => tisd_P3WRDATA_P3CLK(1),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(1),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(1),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(1),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(10),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(10),
          TestSignal => P3WRDATA_P3CLK_dly(10),
          TestSignalName => "P3WRDATA(10)",
          TestDelay => tisd_P3WRDATA_P3CLK(10),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(10),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(10),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(10),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(11),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(11),
          TestSignal => P3WRDATA_P3CLK_dly(11),
          TestSignalName => "P3WRDATA(11)",
          TestDelay => tisd_P3WRDATA_P3CLK(11),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(11),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(11),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(11),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(12),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(12),
          TestSignal => P3WRDATA_P3CLK_dly(12),
          TestSignalName => "P3WRDATA(12)",
          TestDelay => tisd_P3WRDATA_P3CLK(12),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(12),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(12),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(12),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(13),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(13),
          TestSignal => P3WRDATA_P3CLK_dly(13),
          TestSignalName => "P3WRDATA(13)",
          TestDelay => tisd_P3WRDATA_P3CLK(13),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(13),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(13),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(13),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(14),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(14),
          TestSignal => P3WRDATA_P3CLK_dly(14),
          TestSignalName => "P3WRDATA(14)",
          TestDelay => tisd_P3WRDATA_P3CLK(14),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(14),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(14),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(14),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(15),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(15),
          TestSignal => P3WRDATA_P3CLK_dly(15),
          TestSignalName => "P3WRDATA(15)",
          TestDelay => tisd_P3WRDATA_P3CLK(15),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(15),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(15),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(15),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(15),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(16),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(16),
          TestSignal => P3WRDATA_P3CLK_dly(16),
          TestSignalName => "P3WRDATA(16)",
          TestDelay => tisd_P3WRDATA_P3CLK(16),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(16),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(16),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(16),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(16),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(17),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(17),
          TestSignal => P3WRDATA_P3CLK_dly(17),
          TestSignalName => "P3WRDATA(17)",
          TestDelay => tisd_P3WRDATA_P3CLK(17),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(17),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(17),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(17),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(17),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(18),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(18),
          TestSignal => P3WRDATA_P3CLK_dly(18),
          TestSignalName => "P3WRDATA(18)",
          TestDelay => tisd_P3WRDATA_P3CLK(18),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(18),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(18),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(18),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(18),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(19),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(19),
          TestSignal => P3WRDATA_P3CLK_dly(19),
          TestSignalName => "P3WRDATA(19)",
          TestDelay => tisd_P3WRDATA_P3CLK(19),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(19),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(19),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(19),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(19),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(2),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(2),
          TestSignal => P3WRDATA_P3CLK_dly(2),
          TestSignalName => "P3WRDATA(2)",
          TestDelay => tisd_P3WRDATA_P3CLK(2),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(2),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(2),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(2),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(20),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(20),
          TestSignal => P3WRDATA_P3CLK_dly(20),
          TestSignalName => "P3WRDATA(20)",
          TestDelay => tisd_P3WRDATA_P3CLK(20),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(20),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(20),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(20),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(20),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(21),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(21),
          TestSignal => P3WRDATA_P3CLK_dly(21),
          TestSignalName => "P3WRDATA(21)",
          TestDelay => tisd_P3WRDATA_P3CLK(21),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(21),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(21),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(21),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(21),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(22),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(22),
          TestSignal => P3WRDATA_P3CLK_dly(22),
          TestSignalName => "P3WRDATA(22)",
          TestDelay => tisd_P3WRDATA_P3CLK(22),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(22),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(22),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(22),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(22),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(23),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(23),
          TestSignal => P3WRDATA_P3CLK_dly(23),
          TestSignalName => "P3WRDATA(23)",
          TestDelay => tisd_P3WRDATA_P3CLK(23),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(23),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(23),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(23),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(23),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(24),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(24),
          TestSignal => P3WRDATA_P3CLK_dly(24),
          TestSignalName => "P3WRDATA(24)",
          TestDelay => tisd_P3WRDATA_P3CLK(24),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(24),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(24),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(24),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(24),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(25),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(25),
          TestSignal => P3WRDATA_P3CLK_dly(25),
          TestSignalName => "P3WRDATA(25)",
          TestDelay => tisd_P3WRDATA_P3CLK(25),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(25),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(25),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(25),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(25),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(26),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(26),
          TestSignal => P3WRDATA_P3CLK_dly(26),
          TestSignalName => "P3WRDATA(26)",
          TestDelay => tisd_P3WRDATA_P3CLK(26),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(26),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(26),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(26),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(26),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(27),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(27),
          TestSignal => P3WRDATA_P3CLK_dly(27),
          TestSignalName => "P3WRDATA(27)",
          TestDelay => tisd_P3WRDATA_P3CLK(27),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(27),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(27),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(27),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(27),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(28),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(28),
          TestSignal => P3WRDATA_P3CLK_dly(28),
          TestSignalName => "P3WRDATA(28)",
          TestDelay => tisd_P3WRDATA_P3CLK(28),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(28),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(28),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(28),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(28),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(29),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(29),
          TestSignal => P3WRDATA_P3CLK_dly(29),
          TestSignalName => "P3WRDATA(29)",
          TestDelay => tisd_P3WRDATA_P3CLK(29),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(29),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(29),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(29),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(29),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(3),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(3),
          TestSignal => P3WRDATA_P3CLK_dly(3),
          TestSignalName => "P3WRDATA(3)",
          TestDelay => tisd_P3WRDATA_P3CLK(3),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(3),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(3),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(3),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(30),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(30),
          TestSignal => P3WRDATA_P3CLK_dly(30),
          TestSignalName => "P3WRDATA(30)",
          TestDelay => tisd_P3WRDATA_P3CLK(30),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(30),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(30),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(30),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(30),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(31),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(31),
          TestSignal => P3WRDATA_P3CLK_dly(31),
          TestSignalName => "P3WRDATA(31)",
          TestDelay => tisd_P3WRDATA_P3CLK(31),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(31),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(31),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(31),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(31),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(4),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(4),
          TestSignal => P3WRDATA_P3CLK_dly(4),
          TestSignalName => "P3WRDATA(4)",
          TestDelay => tisd_P3WRDATA_P3CLK(4),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(4),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(4),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(4),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(5),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(5),
          TestSignal => P3WRDATA_P3CLK_dly(5),
          TestSignalName => "P3WRDATA(5)",
          TestDelay => tisd_P3WRDATA_P3CLK(5),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(5),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(5),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(5),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(6),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(6),
          TestSignal => P3WRDATA_P3CLK_dly(6),
          TestSignalName => "P3WRDATA(6)",
          TestDelay => tisd_P3WRDATA_P3CLK(6),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(6),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(6),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(6),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(7),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(7),
          TestSignal => P3WRDATA_P3CLK_dly(7),
          TestSignalName => "P3WRDATA(7)",
          TestDelay => tisd_P3WRDATA_P3CLK(7),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(7),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(7),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(7),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(8),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(8),
          TestSignal => P3WRDATA_P3CLK_dly(8),
          TestSignalName => "P3WRDATA(8)",
          TestDelay => tisd_P3WRDATA_P3CLK(8),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(8),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(8),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(8),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRDATA_P3CLK_posedge(9),
          TimingData => Tmkr_P3WRDATA_P3CLK_posedge(9),
          TestSignal => P3WRDATA_P3CLK_dly(9),
          TestSignalName => "P3WRDATA(9)",
          TestDelay => tisd_P3WRDATA_P3CLK(9),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRDATA_P3CLK_posedge_posedge(9),
          HoldHigh => thold_P3WRDATA_P3CLK_posedge_posedge(9),
          SetupLow => tsetup_P3WRDATA_P3CLK_negedge_posedge(9),
          HoldLow => thold_P3WRDATA_P3CLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRMASK_P3CLK_posedge(0),
          TimingData => Tmkr_P3WRMASK_P3CLK_posedge(0),
          TestSignal => P3WRMASK_P3CLK_dly(0),
          TestSignalName => "P3WRMASK(0)",
          TestDelay => tisd_P3WRMASK_P3CLK(0),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRMASK_P3CLK_posedge_posedge(0),
          HoldHigh => thold_P3WRMASK_P3CLK_posedge_posedge(0),
          SetupLow => tsetup_P3WRMASK_P3CLK_negedge_posedge(0),
          HoldLow => thold_P3WRMASK_P3CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRMASK_P3CLK_posedge(1),
          TimingData => Tmkr_P3WRMASK_P3CLK_posedge(1),
          TestSignal => P3WRMASK_P3CLK_dly(1),
          TestSignalName => "P3WRMASK(1)",
          TestDelay => tisd_P3WRMASK_P3CLK(1),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRMASK_P3CLK_posedge_posedge(1),
          HoldHigh => thold_P3WRMASK_P3CLK_posedge_posedge(1),
          SetupLow => tsetup_P3WRMASK_P3CLK_negedge_posedge(1),
          HoldLow => thold_P3WRMASK_P3CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRMASK_P3CLK_posedge(2),
          TimingData => Tmkr_P3WRMASK_P3CLK_posedge(2),
          TestSignal => P3WRMASK_P3CLK_dly(2),
          TestSignalName => "P3WRMASK(2)",
          TestDelay => tisd_P3WRMASK_P3CLK(2),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRMASK_P3CLK_posedge_posedge(2),
          HoldHigh => thold_P3WRMASK_P3CLK_posedge_posedge(2),
          SetupLow => tsetup_P3WRMASK_P3CLK_negedge_posedge(2),
          HoldLow => thold_P3WRMASK_P3CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P3WRMASK_P3CLK_posedge(3),
          TimingData => Tmkr_P3WRMASK_P3CLK_posedge(3),
          TestSignal => P3WRMASK_P3CLK_dly(3),
          TestSignalName => "P3WRMASK(3)",
          TestDelay => tisd_P3WRMASK_P3CLK(3),
          RefSignal => P3CLK_dly,
          RefSignalName => "P3CLK",
          RefDelay => ticd_P3CLK,
          SetupHigh => tsetup_P3WRMASK_P3CLK_posedge_posedge(3),
          HoldHigh => thold_P3WRMASK_P3CLK_posedge_posedge(3),
          SetupLow => tsetup_P3WRMASK_P3CLK_negedge_posedge(3),
          HoldLow => thold_P3WRMASK_P3CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4ARBEN_PLLCLK_posedge(0),
          TimingData => Tmkr_P4ARBEN_PLLCLK_posedge(0),
          TestSignal => P4ARBEN_PLLCLK_dly(0),
          TestSignalName => "P4ARBEN",
          TestDelay => tisd_P4ARBEN_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_P4ARBEN_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_P4ARBEN_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_P4ARBEN_PLLCLK_negedge_posedge(0),
          HoldLow => thold_P4ARBEN_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
         VitalSetupHoldCheck
        (
          Violation => Tviol_P4ARBEN_PLLCLK_posedge(1),
          TimingData => Tmkr_P4ARBEN_PLLCLK_posedge(1),
          TestSignal => P4ARBEN_PLLCLK_dly(1),
          TestSignalName => "P4ARBEN",
          TestDelay => tisd_P4ARBEN_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_P4ARBEN_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_P4ARBEN_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_P4ARBEN_PLLCLK_negedge_posedge(1),
          HoldLow => thold_P4ARBEN_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBA_P4CMDCLK_posedge(0),
          TimingData => Tmkr_P4CMDBA_P4CMDCLK_posedge(0),
          TestSignal => P4CMDBA_P4CMDCLK_dly(0),
          TestSignalName => "P4CMDBA(0)",
          TestDelay => tisd_P4CMDBA_P4CMDCLK(0),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBA_P4CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P4CMDBA_P4CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P4CMDBA_P4CMDCLK_negedge_posedge(0),
          HoldLow => thold_P4CMDBA_P4CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBA_P4CMDCLK_posedge(1),
          TimingData => Tmkr_P4CMDBA_P4CMDCLK_posedge(1),
          TestSignal => P4CMDBA_P4CMDCLK_dly(1),
          TestSignalName => "P4CMDBA(1)",
          TestDelay => tisd_P4CMDBA_P4CMDCLK(1),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBA_P4CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P4CMDBA_P4CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P4CMDBA_P4CMDCLK_negedge_posedge(1),
          HoldLow => thold_P4CMDBA_P4CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBA_P4CMDCLK_posedge(2),
          TimingData => Tmkr_P4CMDBA_P4CMDCLK_posedge(2),
          TestSignal => P4CMDBA_P4CMDCLK_dly(2),
          TestSignalName => "P4CMDBA(2)",
          TestDelay => tisd_P4CMDBA_P4CMDCLK(2),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBA_P4CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P4CMDBA_P4CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P4CMDBA_P4CMDCLK_negedge_posedge(2),
          HoldLow => thold_P4CMDBA_P4CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBL_P4CMDCLK_posedge(0),
          TimingData => Tmkr_P4CMDBL_P4CMDCLK_posedge(0),
          TestSignal => P4CMDBL_P4CMDCLK_dly(0),
          TestSignalName => "P4CMDBL(0)",
          TestDelay => tisd_P4CMDBL_P4CMDCLK(0),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBL_P4CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P4CMDBL_P4CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P4CMDBL_P4CMDCLK_negedge_posedge(0),
          HoldLow => thold_P4CMDBL_P4CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBL_P4CMDCLK_posedge(1),
          TimingData => Tmkr_P4CMDBL_P4CMDCLK_posedge(1),
          TestSignal => P4CMDBL_P4CMDCLK_dly(1),
          TestSignalName => "P4CMDBL(1)",
          TestDelay => tisd_P4CMDBL_P4CMDCLK(1),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBL_P4CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P4CMDBL_P4CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P4CMDBL_P4CMDCLK_negedge_posedge(1),
          HoldLow => thold_P4CMDBL_P4CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBL_P4CMDCLK_posedge(2),
          TimingData => Tmkr_P4CMDBL_P4CMDCLK_posedge(2),
          TestSignal => P4CMDBL_P4CMDCLK_dly(2),
          TestSignalName => "P4CMDBL(2)",
          TestDelay => tisd_P4CMDBL_P4CMDCLK(2),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBL_P4CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P4CMDBL_P4CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P4CMDBL_P4CMDCLK_negedge_posedge(2),
          HoldLow => thold_P4CMDBL_P4CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBL_P4CMDCLK_posedge(3),
          TimingData => Tmkr_P4CMDBL_P4CMDCLK_posedge(3),
          TestSignal => P4CMDBL_P4CMDCLK_dly(3),
          TestSignalName => "P4CMDBL(3)",
          TestDelay => tisd_P4CMDBL_P4CMDCLK(3),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBL_P4CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P4CMDBL_P4CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P4CMDBL_P4CMDCLK_negedge_posedge(3),
          HoldLow => thold_P4CMDBL_P4CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBL_P4CMDCLK_posedge(4),
          TimingData => Tmkr_P4CMDBL_P4CMDCLK_posedge(4),
          TestSignal => P4CMDBL_P4CMDCLK_dly(4),
          TestSignalName => "P4CMDBL(4)",
          TestDelay => tisd_P4CMDBL_P4CMDCLK(4),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBL_P4CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P4CMDBL_P4CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P4CMDBL_P4CMDCLK_negedge_posedge(4),
          HoldLow => thold_P4CMDBL_P4CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDBL_P4CMDCLK_posedge(5),
          TimingData => Tmkr_P4CMDBL_P4CMDCLK_posedge(5),
          TestSignal => P4CMDBL_P4CMDCLK_dly(5),
          TestSignalName => "P4CMDBL(5)",
          TestDelay => tisd_P4CMDBL_P4CMDCLK(5),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDBL_P4CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P4CMDBL_P4CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P4CMDBL_P4CMDCLK_negedge_posedge(5),
          HoldLow => thold_P4CMDBL_P4CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(0),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(0),
          TestSignal => P4CMDCA_P4CMDCLK_dly(0),
          TestSignalName => "P4CMDCA(0)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(0),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(0),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(1),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(1),
          TestSignal => P4CMDCA_P4CMDCLK_dly(1),
          TestSignalName => "P4CMDCA(1)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(1),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(1),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(10),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(10),
          TestSignal => P4CMDCA_P4CMDCLK_dly(10),
          TestSignalName => "P4CMDCA(10)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(10),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(10),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(11),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(11),
          TestSignal => P4CMDCA_P4CMDCLK_dly(11),
          TestSignalName => "P4CMDCA(11)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(11),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(11),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(2),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(2),
          TestSignal => P4CMDCA_P4CMDCLK_dly(2),
          TestSignalName => "P4CMDCA(2)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(2),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(2),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(3),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(3),
          TestSignal => P4CMDCA_P4CMDCLK_dly(3),
          TestSignalName => "P4CMDCA(3)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(3),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(3),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(4),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(4),
          TestSignal => P4CMDCA_P4CMDCLK_dly(4),
          TestSignalName => "P4CMDCA(4)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(4),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(4),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(5),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(5),
          TestSignal => P4CMDCA_P4CMDCLK_dly(5),
          TestSignalName => "P4CMDCA(5)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(5),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(5),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(6),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(6),
          TestSignal => P4CMDCA_P4CMDCLK_dly(6),
          TestSignalName => "P4CMDCA(6)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(6),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(6),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(7),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(7),
          TestSignal => P4CMDCA_P4CMDCLK_dly(7),
          TestSignalName => "P4CMDCA(7)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(7),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(7),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(8),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(8),
          TestSignal => P4CMDCA_P4CMDCLK_dly(8),
          TestSignalName => "P4CMDCA(8)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(8),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(8),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDCA_P4CMDCLK_posedge(9),
          TimingData => Tmkr_P4CMDCA_P4CMDCLK_posedge(9),
          TestSignal => P4CMDCA_P4CMDCLK_dly(9),
          TestSignalName => "P4CMDCA(9)",
          TestDelay => tisd_P4CMDCA_P4CMDCLK(9),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDCA_P4CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P4CMDCA_P4CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P4CMDCA_P4CMDCLK_negedge_posedge(9),
          HoldLow => thold_P4CMDCA_P4CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDEN_P4CMDCLK_posedge,
          TimingData => Tmkr_P4CMDEN_P4CMDCLK_posedge,
          TestSignal => P4CMDEN_P4CMDCLK_dly,
          TestSignalName => "P4CMDEN",
          TestDelay => tisd_P4CMDEN_P4CMDCLK,
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDEN_P4CMDCLK_posedge_posedge,
          HoldHigh => thold_P4CMDEN_P4CMDCLK_posedge_posedge,
          SetupLow => tsetup_P4CMDEN_P4CMDCLK_negedge_posedge,
          HoldLow => thold_P4CMDEN_P4CMDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDINSTR_P4CMDCLK_posedge(0),
          TimingData => Tmkr_P4CMDINSTR_P4CMDCLK_posedge(0),
          TestSignal => P4CMDINSTR_P4CMDCLK_dly(0),
          TestSignalName => "P4CMDINSTR(0)",
          TestDelay => tisd_P4CMDINSTR_P4CMDCLK(0),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDINSTR_P4CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P4CMDINSTR_P4CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P4CMDINSTR_P4CMDCLK_negedge_posedge(0),
          HoldLow => thold_P4CMDINSTR_P4CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDINSTR_P4CMDCLK_posedge(1),
          TimingData => Tmkr_P4CMDINSTR_P4CMDCLK_posedge(1),
          TestSignal => P4CMDINSTR_P4CMDCLK_dly(1),
          TestSignalName => "P4CMDINSTR(1)",
          TestDelay => tisd_P4CMDINSTR_P4CMDCLK(1),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDINSTR_P4CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P4CMDINSTR_P4CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P4CMDINSTR_P4CMDCLK_negedge_posedge(1),
          HoldLow => thold_P4CMDINSTR_P4CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDINSTR_P4CMDCLK_posedge(2),
          TimingData => Tmkr_P4CMDINSTR_P4CMDCLK_posedge(2),
          TestSignal => P4CMDINSTR_P4CMDCLK_dly(2),
          TestSignalName => "P4CMDINSTR(2)",
          TestDelay => tisd_P4CMDINSTR_P4CMDCLK(2),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDINSTR_P4CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P4CMDINSTR_P4CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P4CMDINSTR_P4CMDCLK_negedge_posedge(2),
          HoldLow => thold_P4CMDINSTR_P4CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(0),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(0),
          TestSignal => P4CMDRA_P4CMDCLK_dly(0),
          TestSignalName => "P4CMDRA(0)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(0),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(0),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(1),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(1),
          TestSignal => P4CMDRA_P4CMDCLK_dly(1),
          TestSignalName => "P4CMDRA(1)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(1),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(1),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(10),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(10),
          TestSignal => P4CMDRA_P4CMDCLK_dly(10),
          TestSignalName => "P4CMDRA(10)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(10),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(10),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(11),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(11),
          TestSignal => P4CMDRA_P4CMDCLK_dly(11),
          TestSignalName => "P4CMDRA(11)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(11),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(11),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(12),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(12),
          TestSignal => P4CMDRA_P4CMDCLK_dly(12),
          TestSignalName => "P4CMDRA(12)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(12),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(12),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(12),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(12),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(13),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(13),
          TestSignal => P4CMDRA_P4CMDCLK_dly(13),
          TestSignalName => "P4CMDRA(13)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(13),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(13),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(13),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(13),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(14),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(14),
          TestSignal => P4CMDRA_P4CMDCLK_dly(14),
          TestSignalName => "P4CMDRA(14)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(14),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(14),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(14),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(14),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(2),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(2),
          TestSignal => P4CMDRA_P4CMDCLK_dly(2),
          TestSignalName => "P4CMDRA(2)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(2),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(2),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(3),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(3),
          TestSignal => P4CMDRA_P4CMDCLK_dly(3),
          TestSignalName => "P4CMDRA(3)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(3),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(3),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(4),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(4),
          TestSignal => P4CMDRA_P4CMDCLK_dly(4),
          TestSignalName => "P4CMDRA(4)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(4),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(4),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(5),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(5),
          TestSignal => P4CMDRA_P4CMDCLK_dly(5),
          TestSignalName => "P4CMDRA(5)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(5),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(5),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(6),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(6),
          TestSignal => P4CMDRA_P4CMDCLK_dly(6),
          TestSignalName => "P4CMDRA(6)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(6),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(6),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(7),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(7),
          TestSignal => P4CMDRA_P4CMDCLK_dly(7),
          TestSignalName => "P4CMDRA(7)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(7),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(7),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(8),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(8),
          TestSignal => P4CMDRA_P4CMDCLK_dly(8),
          TestSignalName => "P4CMDRA(8)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(8),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(8),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4CMDRA_P4CMDCLK_posedge(9),
          TimingData => Tmkr_P4CMDRA_P4CMDCLK_posedge(9),
          TestSignal => P4CMDRA_P4CMDCLK_dly(9),
          TestSignalName => "P4CMDRA(9)",
          TestDelay => tisd_P4CMDRA_P4CMDCLK(9),
          RefSignal => P4CMDCLK_dly,
          RefSignalName => "P4CMDCLK",
          RefDelay => ticd_P4CMDCLK,
          SetupHigh => tsetup_P4CMDRA_P4CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P4CMDRA_P4CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P4CMDRA_P4CMDCLK_negedge_posedge(9),
          HoldLow => thold_P4CMDRA_P4CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4EN_P4CLK_posedge,
          TimingData => Tmkr_P4EN_P4CLK_posedge,
          TestSignal => P4EN_P4CLK_dly,
          TestSignalName => "P4EN",
          TestDelay => tisd_P4EN_P4CLK,
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4EN_P4CLK_posedge_posedge,
          HoldHigh => thold_P4EN_P4CLK_posedge_posedge,
          SetupLow => tsetup_P4EN_P4CLK_negedge_posedge,
          HoldLow => thold_P4EN_P4CLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(0),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(0),
          TestSignal => P4WRDATA_P4CLK_dly(0),
          TestSignalName => "P4WRDATA(0)",
          TestDelay => tisd_P4WRDATA_P4CLK(0),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(0),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(0),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(0),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(1),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(1),
          TestSignal => P4WRDATA_P4CLK_dly(1),
          TestSignalName => "P4WRDATA(1)",
          TestDelay => tisd_P4WRDATA_P4CLK(1),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(1),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(1),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(1),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(10),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(10),
          TestSignal => P4WRDATA_P4CLK_dly(10),
          TestSignalName => "P4WRDATA(10)",
          TestDelay => tisd_P4WRDATA_P4CLK(10),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(10),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(10),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(10),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(11),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(11),
          TestSignal => P4WRDATA_P4CLK_dly(11),
          TestSignalName => "P4WRDATA(11)",
          TestDelay => tisd_P4WRDATA_P4CLK(11),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(11),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(11),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(11),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(12),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(12),
          TestSignal => P4WRDATA_P4CLK_dly(12),
          TestSignalName => "P4WRDATA(12)",
          TestDelay => tisd_P4WRDATA_P4CLK(12),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(12),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(12),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(12),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(13),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(13),
          TestSignal => P4WRDATA_P4CLK_dly(13),
          TestSignalName => "P4WRDATA(13)",
          TestDelay => tisd_P4WRDATA_P4CLK(13),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(13),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(13),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(13),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(14),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(14),
          TestSignal => P4WRDATA_P4CLK_dly(14),
          TestSignalName => "P4WRDATA(14)",
          TestDelay => tisd_P4WRDATA_P4CLK(14),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(14),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(14),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(14),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(15),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(15),
          TestSignal => P4WRDATA_P4CLK_dly(15),
          TestSignalName => "P4WRDATA(15)",
          TestDelay => tisd_P4WRDATA_P4CLK(15),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(15),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(15),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(15),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(15),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(16),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(16),
          TestSignal => P4WRDATA_P4CLK_dly(16),
          TestSignalName => "P4WRDATA(16)",
          TestDelay => tisd_P4WRDATA_P4CLK(16),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(16),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(16),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(16),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(16),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(17),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(17),
          TestSignal => P4WRDATA_P4CLK_dly(17),
          TestSignalName => "P4WRDATA(17)",
          TestDelay => tisd_P4WRDATA_P4CLK(17),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(17),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(17),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(17),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(17),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(18),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(18),
          TestSignal => P4WRDATA_P4CLK_dly(18),
          TestSignalName => "P4WRDATA(18)",
          TestDelay => tisd_P4WRDATA_P4CLK(18),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(18),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(18),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(18),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(18),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(19),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(19),
          TestSignal => P4WRDATA_P4CLK_dly(19),
          TestSignalName => "P4WRDATA(19)",
          TestDelay => tisd_P4WRDATA_P4CLK(19),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(19),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(19),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(19),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(19),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(2),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(2),
          TestSignal => P4WRDATA_P4CLK_dly(2),
          TestSignalName => "P4WRDATA(2)",
          TestDelay => tisd_P4WRDATA_P4CLK(2),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(2),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(2),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(2),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(20),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(20),
          TestSignal => P4WRDATA_P4CLK_dly(20),
          TestSignalName => "P4WRDATA(20)",
          TestDelay => tisd_P4WRDATA_P4CLK(20),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(20),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(20),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(20),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(20),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(21),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(21),
          TestSignal => P4WRDATA_P4CLK_dly(21),
          TestSignalName => "P4WRDATA(21)",
          TestDelay => tisd_P4WRDATA_P4CLK(21),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(21),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(21),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(21),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(21),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(22),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(22),
          TestSignal => P4WRDATA_P4CLK_dly(22),
          TestSignalName => "P4WRDATA(22)",
          TestDelay => tisd_P4WRDATA_P4CLK(22),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(22),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(22),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(22),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(22),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(23),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(23),
          TestSignal => P4WRDATA_P4CLK_dly(23),
          TestSignalName => "P4WRDATA(23)",
          TestDelay => tisd_P4WRDATA_P4CLK(23),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(23),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(23),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(23),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(23),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(24),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(24),
          TestSignal => P4WRDATA_P4CLK_dly(24),
          TestSignalName => "P4WRDATA(24)",
          TestDelay => tisd_P4WRDATA_P4CLK(24),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(24),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(24),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(24),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(24),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(25),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(25),
          TestSignal => P4WRDATA_P4CLK_dly(25),
          TestSignalName => "P4WRDATA(25)",
          TestDelay => tisd_P4WRDATA_P4CLK(25),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(25),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(25),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(25),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(25),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(26),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(26),
          TestSignal => P4WRDATA_P4CLK_dly(26),
          TestSignalName => "P4WRDATA(26)",
          TestDelay => tisd_P4WRDATA_P4CLK(26),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(26),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(26),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(26),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(26),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(27),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(27),
          TestSignal => P4WRDATA_P4CLK_dly(27),
          TestSignalName => "P4WRDATA(27)",
          TestDelay => tisd_P4WRDATA_P4CLK(27),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(27),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(27),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(27),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(27),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(28),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(28),
          TestSignal => P4WRDATA_P4CLK_dly(28),
          TestSignalName => "P4WRDATA(28)",
          TestDelay => tisd_P4WRDATA_P4CLK(28),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(28),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(28),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(28),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(28),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(29),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(29),
          TestSignal => P4WRDATA_P4CLK_dly(29),
          TestSignalName => "P4WRDATA(29)",
          TestDelay => tisd_P4WRDATA_P4CLK(29),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(29),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(29),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(29),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(29),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(3),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(3),
          TestSignal => P4WRDATA_P4CLK_dly(3),
          TestSignalName => "P4WRDATA(3)",
          TestDelay => tisd_P4WRDATA_P4CLK(3),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(3),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(3),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(3),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(30),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(30),
          TestSignal => P4WRDATA_P4CLK_dly(30),
          TestSignalName => "P4WRDATA(30)",
          TestDelay => tisd_P4WRDATA_P4CLK(30),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(30),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(30),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(30),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(30),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(31),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(31),
          TestSignal => P4WRDATA_P4CLK_dly(31),
          TestSignalName => "P4WRDATA(31)",
          TestDelay => tisd_P4WRDATA_P4CLK(31),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(31),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(31),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(31),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(31),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(4),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(4),
          TestSignal => P4WRDATA_P4CLK_dly(4),
          TestSignalName => "P4WRDATA(4)",
          TestDelay => tisd_P4WRDATA_P4CLK(4),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(4),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(4),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(4),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(5),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(5),
          TestSignal => P4WRDATA_P4CLK_dly(5),
          TestSignalName => "P4WRDATA(5)",
          TestDelay => tisd_P4WRDATA_P4CLK(5),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(5),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(5),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(5),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(6),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(6),
          TestSignal => P4WRDATA_P4CLK_dly(6),
          TestSignalName => "P4WRDATA(6)",
          TestDelay => tisd_P4WRDATA_P4CLK(6),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(6),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(6),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(6),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(7),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(7),
          TestSignal => P4WRDATA_P4CLK_dly(7),
          TestSignalName => "P4WRDATA(7)",
          TestDelay => tisd_P4WRDATA_P4CLK(7),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(7),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(7),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(7),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(8),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(8),
          TestSignal => P4WRDATA_P4CLK_dly(8),
          TestSignalName => "P4WRDATA(8)",
          TestDelay => tisd_P4WRDATA_P4CLK(8),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(8),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(8),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(8),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRDATA_P4CLK_posedge(9),
          TimingData => Tmkr_P4WRDATA_P4CLK_posedge(9),
          TestSignal => P4WRDATA_P4CLK_dly(9),
          TestSignalName => "P4WRDATA(9)",
          TestDelay => tisd_P4WRDATA_P4CLK(9),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRDATA_P4CLK_posedge_posedge(9),
          HoldHigh => thold_P4WRDATA_P4CLK_posedge_posedge(9),
          SetupLow => tsetup_P4WRDATA_P4CLK_negedge_posedge(9),
          HoldLow => thold_P4WRDATA_P4CLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRMASK_P4CLK_posedge(0),
          TimingData => Tmkr_P4WRMASK_P4CLK_posedge(0),
          TestSignal => P4WRMASK_P4CLK_dly(0),
          TestSignalName => "P4WRMASK(0)",
          TestDelay => tisd_P4WRMASK_P4CLK(0),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRMASK_P4CLK_posedge_posedge(0),
          HoldHigh => thold_P4WRMASK_P4CLK_posedge_posedge(0),
          SetupLow => tsetup_P4WRMASK_P4CLK_negedge_posedge(0),
          HoldLow => thold_P4WRMASK_P4CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRMASK_P4CLK_posedge(1),
          TimingData => Tmkr_P4WRMASK_P4CLK_posedge(1),
          TestSignal => P4WRMASK_P4CLK_dly(1),
          TestSignalName => "P4WRMASK(1)",
          TestDelay => tisd_P4WRMASK_P4CLK(1),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRMASK_P4CLK_posedge_posedge(1),
          HoldHigh => thold_P4WRMASK_P4CLK_posedge_posedge(1),
          SetupLow => tsetup_P4WRMASK_P4CLK_negedge_posedge(1),
          HoldLow => thold_P4WRMASK_P4CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRMASK_P4CLK_posedge(2),
          TimingData => Tmkr_P4WRMASK_P4CLK_posedge(2),
          TestSignal => P4WRMASK_P4CLK_dly(2),
          TestSignalName => "P4WRMASK(2)",
          TestDelay => tisd_P4WRMASK_P4CLK(2),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRMASK_P4CLK_posedge_posedge(2),
          HoldHigh => thold_P4WRMASK_P4CLK_posedge_posedge(2),
          SetupLow => tsetup_P4WRMASK_P4CLK_negedge_posedge(2),
          HoldLow => thold_P4WRMASK_P4CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P4WRMASK_P4CLK_posedge(3),
          TimingData => Tmkr_P4WRMASK_P4CLK_posedge(3),
          TestSignal => P4WRMASK_P4CLK_dly(3),
          TestSignalName => "P4WRMASK(3)",
          TestDelay => tisd_P4WRMASK_P4CLK(3),
          RefSignal => P4CLK_dly,
          RefSignalName => "P4CLK",
          RefDelay => ticd_P4CLK,
          SetupHigh => tsetup_P4WRMASK_P4CLK_posedge_posedge(3),
          HoldHigh => thold_P4WRMASK_P4CLK_posedge_posedge(3),
          SetupLow => tsetup_P4WRMASK_P4CLK_negedge_posedge(3),
          HoldLow => thold_P4WRMASK_P4CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5ARBEN_PLLCLK_posedge(0),
          TimingData => Tmkr_P5ARBEN_PLLCLK_posedge(0),
          TestSignal => P5ARBEN_PLLCLK_dly(0),
          TestSignalName => "P5ARBEN",
          TestDelay => tisd_P5ARBEN_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_P5ARBEN_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_P5ARBEN_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_P5ARBEN_PLLCLK_negedge_posedge(0),
          HoldLow => thold_P5ARBEN_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5ARBEN_PLLCLK_posedge(1),
          TimingData => Tmkr_P5ARBEN_PLLCLK_posedge(1),
          TestSignal => P5ARBEN_PLLCLK_dly(1),
          TestSignalName => "P5ARBEN",
          TestDelay => tisd_P5ARBEN_PLLCLK(1),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_P5ARBEN_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_P5ARBEN_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_P5ARBEN_PLLCLK_negedge_posedge(1),
          HoldLow => thold_P5ARBEN_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBA_P5CMDCLK_posedge(0),
          TimingData => Tmkr_P5CMDBA_P5CMDCLK_posedge(0),
          TestSignal => P5CMDBA_P5CMDCLK_dly(0),
          TestSignalName => "P5CMDBA(0)",
          TestDelay => tisd_P5CMDBA_P5CMDCLK(0),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBA_P5CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P5CMDBA_P5CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P5CMDBA_P5CMDCLK_negedge_posedge(0),
          HoldLow => thold_P5CMDBA_P5CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBA_P5CMDCLK_posedge(1),
          TimingData => Tmkr_P5CMDBA_P5CMDCLK_posedge(1),
          TestSignal => P5CMDBA_P5CMDCLK_dly(1),
          TestSignalName => "P5CMDBA(1)",
          TestDelay => tisd_P5CMDBA_P5CMDCLK(1),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBA_P5CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P5CMDBA_P5CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P5CMDBA_P5CMDCLK_negedge_posedge(1),
          HoldLow => thold_P5CMDBA_P5CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBA_P5CMDCLK_posedge(2),
          TimingData => Tmkr_P5CMDBA_P5CMDCLK_posedge(2),
          TestSignal => P5CMDBA_P5CMDCLK_dly(2),
          TestSignalName => "P5CMDBA(2)",
          TestDelay => tisd_P5CMDBA_P5CMDCLK(2),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBA_P5CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P5CMDBA_P5CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P5CMDBA_P5CMDCLK_negedge_posedge(2),
          HoldLow => thold_P5CMDBA_P5CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBL_P5CMDCLK_posedge(0),
          TimingData => Tmkr_P5CMDBL_P5CMDCLK_posedge(0),
          TestSignal => P5CMDBL_P5CMDCLK_dly(0),
          TestSignalName => "P5CMDBL(0)",
          TestDelay => tisd_P5CMDBL_P5CMDCLK(0),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBL_P5CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P5CMDBL_P5CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P5CMDBL_P5CMDCLK_negedge_posedge(0),
          HoldLow => thold_P5CMDBL_P5CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBL_P5CMDCLK_posedge(1),
          TimingData => Tmkr_P5CMDBL_P5CMDCLK_posedge(1),
          TestSignal => P5CMDBL_P5CMDCLK_dly(1),
          TestSignalName => "P5CMDBL(1)",
          TestDelay => tisd_P5CMDBL_P5CMDCLK(1),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBL_P5CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P5CMDBL_P5CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P5CMDBL_P5CMDCLK_negedge_posedge(1),
          HoldLow => thold_P5CMDBL_P5CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBL_P5CMDCLK_posedge(2),
          TimingData => Tmkr_P5CMDBL_P5CMDCLK_posedge(2),
          TestSignal => P5CMDBL_P5CMDCLK_dly(2),
          TestSignalName => "P5CMDBL(2)",
          TestDelay => tisd_P5CMDBL_P5CMDCLK(2),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBL_P5CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P5CMDBL_P5CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P5CMDBL_P5CMDCLK_negedge_posedge(2),
          HoldLow => thold_P5CMDBL_P5CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBL_P5CMDCLK_posedge(3),
          TimingData => Tmkr_P5CMDBL_P5CMDCLK_posedge(3),
          TestSignal => P5CMDBL_P5CMDCLK_dly(3),
          TestSignalName => "P5CMDBL(3)",
          TestDelay => tisd_P5CMDBL_P5CMDCLK(3),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBL_P5CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P5CMDBL_P5CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P5CMDBL_P5CMDCLK_negedge_posedge(3),
          HoldLow => thold_P5CMDBL_P5CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBL_P5CMDCLK_posedge(4),
          TimingData => Tmkr_P5CMDBL_P5CMDCLK_posedge(4),
          TestSignal => P5CMDBL_P5CMDCLK_dly(4),
          TestSignalName => "P5CMDBL(4)",
          TestDelay => tisd_P5CMDBL_P5CMDCLK(4),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBL_P5CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P5CMDBL_P5CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P5CMDBL_P5CMDCLK_negedge_posedge(4),
          HoldLow => thold_P5CMDBL_P5CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDBL_P5CMDCLK_posedge(5),
          TimingData => Tmkr_P5CMDBL_P5CMDCLK_posedge(5),
          TestSignal => P5CMDBL_P5CMDCLK_dly(5),
          TestSignalName => "P5CMDBL(5)",
          TestDelay => tisd_P5CMDBL_P5CMDCLK(5),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDBL_P5CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P5CMDBL_P5CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P5CMDBL_P5CMDCLK_negedge_posedge(5),
          HoldLow => thold_P5CMDBL_P5CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(0),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(0),
          TestSignal => P5CMDCA_P5CMDCLK_dly(0),
          TestSignalName => "P5CMDCA(0)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(0),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(0),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(1),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(1),
          TestSignal => P5CMDCA_P5CMDCLK_dly(1),
          TestSignalName => "P5CMDCA(1)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(1),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(1),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(10),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(10),
          TestSignal => P5CMDCA_P5CMDCLK_dly(10),
          TestSignalName => "P5CMDCA(10)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(10),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(10),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(11),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(11),
          TestSignal => P5CMDCA_P5CMDCLK_dly(11),
          TestSignalName => "P5CMDCA(11)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(11),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(11),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(2),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(2),
          TestSignal => P5CMDCA_P5CMDCLK_dly(2),
          TestSignalName => "P5CMDCA(2)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(2),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(2),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(3),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(3),
          TestSignal => P5CMDCA_P5CMDCLK_dly(3),
          TestSignalName => "P5CMDCA(3)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(3),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(3),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(4),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(4),
          TestSignal => P5CMDCA_P5CMDCLK_dly(4),
          TestSignalName => "P5CMDCA(4)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(4),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(4),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(5),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(5),
          TestSignal => P5CMDCA_P5CMDCLK_dly(5),
          TestSignalName => "P5CMDCA(5)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(5),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(5),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(6),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(6),
          TestSignal => P5CMDCA_P5CMDCLK_dly(6),
          TestSignalName => "P5CMDCA(6)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(6),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(6),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(7),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(7),
          TestSignal => P5CMDCA_P5CMDCLK_dly(7),
          TestSignalName => "P5CMDCA(7)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(7),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(7),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(8),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(8),
          TestSignal => P5CMDCA_P5CMDCLK_dly(8),
          TestSignalName => "P5CMDCA(8)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(8),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(8),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDCA_P5CMDCLK_posedge(9),
          TimingData => Tmkr_P5CMDCA_P5CMDCLK_posedge(9),
          TestSignal => P5CMDCA_P5CMDCLK_dly(9),
          TestSignalName => "P5CMDCA(9)",
          TestDelay => tisd_P5CMDCA_P5CMDCLK(9),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDCA_P5CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P5CMDCA_P5CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P5CMDCA_P5CMDCLK_negedge_posedge(9),
          HoldLow => thold_P5CMDCA_P5CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDEN_P5CMDCLK_posedge,
          TimingData => Tmkr_P5CMDEN_P5CMDCLK_posedge,
          TestSignal => P5CMDEN_P5CMDCLK_dly,
          TestSignalName => "P5CMDEN",
          TestDelay => tisd_P5CMDEN_P5CMDCLK,
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDEN_P5CMDCLK_posedge_posedge,
          HoldHigh => thold_P5CMDEN_P5CMDCLK_posedge_posedge,
          SetupLow => tsetup_P5CMDEN_P5CMDCLK_negedge_posedge,
          HoldLow => thold_P5CMDEN_P5CMDCLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDINSTR_P5CMDCLK_posedge(0),
          TimingData => Tmkr_P5CMDINSTR_P5CMDCLK_posedge(0),
          TestSignal => P5CMDINSTR_P5CMDCLK_dly(0),
          TestSignalName => "P5CMDINSTR(0)",
          TestDelay => tisd_P5CMDINSTR_P5CMDCLK(0),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDINSTR_P5CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P5CMDINSTR_P5CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P5CMDINSTR_P5CMDCLK_negedge_posedge(0),
          HoldLow => thold_P5CMDINSTR_P5CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDINSTR_P5CMDCLK_posedge(1),
          TimingData => Tmkr_P5CMDINSTR_P5CMDCLK_posedge(1),
          TestSignal => P5CMDINSTR_P5CMDCLK_dly(1),
          TestSignalName => "P5CMDINSTR(1)",
          TestDelay => tisd_P5CMDINSTR_P5CMDCLK(1),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDINSTR_P5CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P5CMDINSTR_P5CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P5CMDINSTR_P5CMDCLK_negedge_posedge(1),
          HoldLow => thold_P5CMDINSTR_P5CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDINSTR_P5CMDCLK_posedge(2),
          TimingData => Tmkr_P5CMDINSTR_P5CMDCLK_posedge(2),
          TestSignal => P5CMDINSTR_P5CMDCLK_dly(2),
          TestSignalName => "P5CMDINSTR(2)",
          TestDelay => tisd_P5CMDINSTR_P5CMDCLK(2),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDINSTR_P5CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P5CMDINSTR_P5CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P5CMDINSTR_P5CMDCLK_negedge_posedge(2),
          HoldLow => thold_P5CMDINSTR_P5CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(0),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(0),
          TestSignal => P5CMDRA_P5CMDCLK_dly(0),
          TestSignalName => "P5CMDRA(0)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(0),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(0),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(0),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(0),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(1),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(1),
          TestSignal => P5CMDRA_P5CMDCLK_dly(1),
          TestSignalName => "P5CMDRA(1)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(1),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(1),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(1),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(1),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(10),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(10),
          TestSignal => P5CMDRA_P5CMDCLK_dly(10),
          TestSignalName => "P5CMDRA(10)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(10),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(10),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(10),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(10),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(11),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(11),
          TestSignal => P5CMDRA_P5CMDCLK_dly(11),
          TestSignalName => "P5CMDRA(11)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(11),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(11),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(11),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(11),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(12),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(12),
          TestSignal => P5CMDRA_P5CMDCLK_dly(12),
          TestSignalName => "P5CMDRA(12)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(12),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(12),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(12),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(12),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(13),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(13),
          TestSignal => P5CMDRA_P5CMDCLK_dly(13),
          TestSignalName => "P5CMDRA(13)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(13),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(13),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(13),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(13),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(14),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(14),
          TestSignal => P5CMDRA_P5CMDCLK_dly(14),
          TestSignalName => "P5CMDRA(14)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(14),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(14),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(14),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(14),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(2),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(2),
          TestSignal => P5CMDRA_P5CMDCLK_dly(2),
          TestSignalName => "P5CMDRA(2)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(2),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(2),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(2),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(2),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(3),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(3),
          TestSignal => P5CMDRA_P5CMDCLK_dly(3),
          TestSignalName => "P5CMDRA(3)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(3),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(3),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(3),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(3),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(4),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(4),
          TestSignal => P5CMDRA_P5CMDCLK_dly(4),
          TestSignalName => "P5CMDRA(4)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(4),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(4),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(4),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(4),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(5),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(5),
          TestSignal => P5CMDRA_P5CMDCLK_dly(5),
          TestSignalName => "P5CMDRA(5)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(5),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(5),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(5),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(5),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(6),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(6),
          TestSignal => P5CMDRA_P5CMDCLK_dly(6),
          TestSignalName => "P5CMDRA(6)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(6),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(6),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(6),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(6),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(7),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(7),
          TestSignal => P5CMDRA_P5CMDCLK_dly(7),
          TestSignalName => "P5CMDRA(7)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(7),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(7),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(7),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(7),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(8),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(8),
          TestSignal => P5CMDRA_P5CMDCLK_dly(8),
          TestSignalName => "P5CMDRA(8)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(8),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(8),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(8),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(8),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5CMDRA_P5CMDCLK_posedge(9),
          TimingData => Tmkr_P5CMDRA_P5CMDCLK_posedge(9),
          TestSignal => P5CMDRA_P5CMDCLK_dly(9),
          TestSignalName => "P5CMDRA(9)",
          TestDelay => tisd_P5CMDRA_P5CMDCLK(9),
          RefSignal => P5CMDCLK_dly,
          RefSignalName => "P5CMDCLK",
          RefDelay => ticd_P5CMDCLK,
          SetupHigh => tsetup_P5CMDRA_P5CMDCLK_posedge_posedge(9),
          HoldHigh => thold_P5CMDRA_P5CMDCLK_posedge_posedge(9),
          SetupLow => tsetup_P5CMDRA_P5CMDCLK_negedge_posedge(9),
          HoldLow => thold_P5CMDRA_P5CMDCLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5EN_P5CLK_posedge,
          TimingData => Tmkr_P5EN_P5CLK_posedge,
          TestSignal => P5EN_P5CLK_dly,
          TestSignalName => "P5EN",
          TestDelay => tisd_P5EN_P5CLK,
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5EN_P5CLK_posedge_posedge,
          HoldHigh => thold_P5EN_P5CLK_posedge_posedge,
          SetupLow => tsetup_P5EN_P5CLK_negedge_posedge,
          HoldLow => thold_P5EN_P5CLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(0),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(0),
          TestSignal => P5WRDATA_P5CLK_dly(0),
          TestSignalName => "P5WRDATA(0)",
          TestDelay => tisd_P5WRDATA_P5CLK(0),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(0),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(0),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(0),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(1),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(1),
          TestSignal => P5WRDATA_P5CLK_dly(1),
          TestSignalName => "P5WRDATA(1)",
          TestDelay => tisd_P5WRDATA_P5CLK(1),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(1),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(1),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(1),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(10),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(10),
          TestSignal => P5WRDATA_P5CLK_dly(10),
          TestSignalName => "P5WRDATA(10)",
          TestDelay => tisd_P5WRDATA_P5CLK(10),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(10),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(10),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(10),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(10),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(11),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(11),
          TestSignal => P5WRDATA_P5CLK_dly(11),
          TestSignalName => "P5WRDATA(11)",
          TestDelay => tisd_P5WRDATA_P5CLK(11),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(11),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(11),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(11),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(11),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(12),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(12),
          TestSignal => P5WRDATA_P5CLK_dly(12),
          TestSignalName => "P5WRDATA(12)",
          TestDelay => tisd_P5WRDATA_P5CLK(12),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(12),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(12),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(12),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(12),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(13),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(13),
          TestSignal => P5WRDATA_P5CLK_dly(13),
          TestSignalName => "P5WRDATA(13)",
          TestDelay => tisd_P5WRDATA_P5CLK(13),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(13),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(13),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(13),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(13),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(14),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(14),
          TestSignal => P5WRDATA_P5CLK_dly(14),
          TestSignalName => "P5WRDATA(14)",
          TestDelay => tisd_P5WRDATA_P5CLK(14),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(14),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(14),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(14),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(14),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(15),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(15),
          TestSignal => P5WRDATA_P5CLK_dly(15),
          TestSignalName => "P5WRDATA(15)",
          TestDelay => tisd_P5WRDATA_P5CLK(15),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(15),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(15),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(15),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(15),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(16),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(16),
          TestSignal => P5WRDATA_P5CLK_dly(16),
          TestSignalName => "P5WRDATA(16)",
          TestDelay => tisd_P5WRDATA_P5CLK(16),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(16),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(16),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(16),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(16),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(17),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(17),
          TestSignal => P5WRDATA_P5CLK_dly(17),
          TestSignalName => "P5WRDATA(17)",
          TestDelay => tisd_P5WRDATA_P5CLK(17),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(17),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(17),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(17),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(17),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(18),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(18),
          TestSignal => P5WRDATA_P5CLK_dly(18),
          TestSignalName => "P5WRDATA(18)",
          TestDelay => tisd_P5WRDATA_P5CLK(18),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(18),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(18),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(18),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(18),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(19),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(19),
          TestSignal => P5WRDATA_P5CLK_dly(19),
          TestSignalName => "P5WRDATA(19)",
          TestDelay => tisd_P5WRDATA_P5CLK(19),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(19),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(19),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(19),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(19),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(2),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(2),
          TestSignal => P5WRDATA_P5CLK_dly(2),
          TestSignalName => "P5WRDATA(2)",
          TestDelay => tisd_P5WRDATA_P5CLK(2),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(2),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(2),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(2),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(20),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(20),
          TestSignal => P5WRDATA_P5CLK_dly(20),
          TestSignalName => "P5WRDATA(20)",
          TestDelay => tisd_P5WRDATA_P5CLK(20),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(20),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(20),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(20),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(20),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(21),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(21),
          TestSignal => P5WRDATA_P5CLK_dly(21),
          TestSignalName => "P5WRDATA(21)",
          TestDelay => tisd_P5WRDATA_P5CLK(21),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(21),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(21),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(21),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(21),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(22),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(22),
          TestSignal => P5WRDATA_P5CLK_dly(22),
          TestSignalName => "P5WRDATA(22)",
          TestDelay => tisd_P5WRDATA_P5CLK(22),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(22),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(22),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(22),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(22),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(23),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(23),
          TestSignal => P5WRDATA_P5CLK_dly(23),
          TestSignalName => "P5WRDATA(23)",
          TestDelay => tisd_P5WRDATA_P5CLK(23),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(23),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(23),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(23),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(23),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(24),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(24),
          TestSignal => P5WRDATA_P5CLK_dly(24),
          TestSignalName => "P5WRDATA(24)",
          TestDelay => tisd_P5WRDATA_P5CLK(24),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(24),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(24),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(24),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(24),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(25),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(25),
          TestSignal => P5WRDATA_P5CLK_dly(25),
          TestSignalName => "P5WRDATA(25)",
          TestDelay => tisd_P5WRDATA_P5CLK(25),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(25),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(25),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(25),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(25),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(26),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(26),
          TestSignal => P5WRDATA_P5CLK_dly(26),
          TestSignalName => "P5WRDATA(26)",
          TestDelay => tisd_P5WRDATA_P5CLK(26),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(26),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(26),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(26),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(26),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(27),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(27),
          TestSignal => P5WRDATA_P5CLK_dly(27),
          TestSignalName => "P5WRDATA(27)",
          TestDelay => tisd_P5WRDATA_P5CLK(27),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(27),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(27),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(27),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(27),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(28),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(28),
          TestSignal => P5WRDATA_P5CLK_dly(28),
          TestSignalName => "P5WRDATA(28)",
          TestDelay => tisd_P5WRDATA_P5CLK(28),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(28),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(28),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(28),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(28),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(29),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(29),
          TestSignal => P5WRDATA_P5CLK_dly(29),
          TestSignalName => "P5WRDATA(29)",
          TestDelay => tisd_P5WRDATA_P5CLK(29),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(29),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(29),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(29),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(29),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(3),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(3),
          TestSignal => P5WRDATA_P5CLK_dly(3),
          TestSignalName => "P5WRDATA(3)",
          TestDelay => tisd_P5WRDATA_P5CLK(3),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(3),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(3),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(3),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(30),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(30),
          TestSignal => P5WRDATA_P5CLK_dly(30),
          TestSignalName => "P5WRDATA(30)",
          TestDelay => tisd_P5WRDATA_P5CLK(30),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(30),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(30),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(30),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(30),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(31),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(31),
          TestSignal => P5WRDATA_P5CLK_dly(31),
          TestSignalName => "P5WRDATA(31)",
          TestDelay => tisd_P5WRDATA_P5CLK(31),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(31),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(31),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(31),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(31),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(4),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(4),
          TestSignal => P5WRDATA_P5CLK_dly(4),
          TestSignalName => "P5WRDATA(4)",
          TestDelay => tisd_P5WRDATA_P5CLK(4),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(4),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(4),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(4),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(5),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(5),
          TestSignal => P5WRDATA_P5CLK_dly(5),
          TestSignalName => "P5WRDATA(5)",
          TestDelay => tisd_P5WRDATA_P5CLK(5),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(5),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(5),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(5),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(5),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(6),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(6),
          TestSignal => P5WRDATA_P5CLK_dly(6),
          TestSignalName => "P5WRDATA(6)",
          TestDelay => tisd_P5WRDATA_P5CLK(6),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(6),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(6),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(6),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(6),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(7),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(7),
          TestSignal => P5WRDATA_P5CLK_dly(7),
          TestSignalName => "P5WRDATA(7)",
          TestDelay => tisd_P5WRDATA_P5CLK(7),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(7),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(7),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(7),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(7),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(8),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(8),
          TestSignal => P5WRDATA_P5CLK_dly(8),
          TestSignalName => "P5WRDATA(8)",
          TestDelay => tisd_P5WRDATA_P5CLK(8),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(8),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(8),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(8),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(8),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRDATA_P5CLK_posedge(9),
          TimingData => Tmkr_P5WRDATA_P5CLK_posedge(9),
          TestSignal => P5WRDATA_P5CLK_dly(9),
          TestSignalName => "P5WRDATA(9)",
          TestDelay => tisd_P5WRDATA_P5CLK(9),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRDATA_P5CLK_posedge_posedge(9),
          HoldHigh => thold_P5WRDATA_P5CLK_posedge_posedge(9),
          SetupLow => tsetup_P5WRDATA_P5CLK_negedge_posedge(9),
          HoldLow => thold_P5WRDATA_P5CLK_negedge_posedge(9),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRMASK_P5CLK_posedge(0),
          TimingData => Tmkr_P5WRMASK_P5CLK_posedge(0),
          TestSignal => P5WRMASK_P5CLK_dly(0),
          TestSignalName => "P5WRMASK(0)",
          TestDelay => tisd_P5WRMASK_P5CLK(0),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRMASK_P5CLK_posedge_posedge(0),
          HoldHigh => thold_P5WRMASK_P5CLK_posedge_posedge(0),
          SetupLow => tsetup_P5WRMASK_P5CLK_negedge_posedge(0),
          HoldLow => thold_P5WRMASK_P5CLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRMASK_P5CLK_posedge(1),
          TimingData => Tmkr_P5WRMASK_P5CLK_posedge(1),
          TestSignal => P5WRMASK_P5CLK_dly(1),
          TestSignalName => "P5WRMASK(1)",
          TestDelay => tisd_P5WRMASK_P5CLK(1),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRMASK_P5CLK_posedge_posedge(1),
          HoldHigh => thold_P5WRMASK_P5CLK_posedge_posedge(1),
          SetupLow => tsetup_P5WRMASK_P5CLK_negedge_posedge(1),
          HoldLow => thold_P5WRMASK_P5CLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRMASK_P5CLK_posedge(2),
          TimingData => Tmkr_P5WRMASK_P5CLK_posedge(2),
          TestSignal => P5WRMASK_P5CLK_dly(2),
          TestSignalName => "P5WRMASK(2)",
          TestDelay => tisd_P5WRMASK_P5CLK(2),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRMASK_P5CLK_posedge_posedge(2),
          HoldHigh => thold_P5WRMASK_P5CLK_posedge_posedge(2),
          SetupLow => tsetup_P5WRMASK_P5CLK_negedge_posedge(2),
          HoldLow => thold_P5WRMASK_P5CLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_P5WRMASK_P5CLK_posedge(3),
          TimingData => Tmkr_P5WRMASK_P5CLK_posedge(3),
          TestSignal => P5WRMASK_P5CLK_dly(3),
          TestSignalName => "P5WRMASK(3)",
          TestDelay => tisd_P5WRMASK_P5CLK(3),
          RefSignal => P5CLK_dly,
          RefSignalName => "P5CLK",
          RefDelay => ticd_P5CLK,
          SetupHigh => tsetup_P5WRMASK_P5CLK_posedge_posedge(3),
          HoldHigh => thold_P5WRMASK_P5CLK_posedge_posedge(3),
          SetupLow => tsetup_P5WRMASK_P5CLK_negedge_posedge(3),
          HoldLow => thold_P5WRMASK_P5CLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_PLLCE_PLLCLK_posedge(0),
          TimingData => Tmkr_PLLCE_PLLCLK_posedge(0),
          TestSignal => PLLCE_PLLCLK_dly(0),
          TestSignalName => "PLLCE(0)",
          TestDelay => tisd_PLLCE_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_PLLCE_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_PLLCE_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_PLLCE_PLLCLK_negedge_posedge(0),
          HoldLow => thold_PLLCE_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_PLLCE_PLLCLK_posedge(1),
          TimingData => Tmkr_PLLCE_PLLCLK_posedge(1),
          TestSignal => PLLCE_PLLCLK_dly(1),
          TestSignalName => "PLLCE(1)",
          TestDelay => tisd_PLLCE_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_PLLCE_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_PLLCE_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_PLLCE_PLLCLK_negedge_posedge(1),
          HoldLow => thold_PLLCE_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_PLLCE_PLLCLK_posedge(2),
          TimingData => Tmkr_PLLCE_PLLCLK_posedge(2),
          TestSignal => PLLCE_PLLCLK_dly(2),
          TestSignalName => "PLLCE(0)",
          TestDelay => tisd_PLLCE_PLLCLK(2),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_PLLCE_PLLCLK_posedge_posedge(2),
          HoldHigh => thold_PLLCE_PLLCLK_posedge_posedge(2),
          SetupLow => tsetup_PLLCE_PLLCLK_negedge_posedge(2),
          HoldLow => thold_PLLCE_PLLCLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_PLLCE_PLLCLK_posedge(3),
          TimingData => Tmkr_PLLCE_PLLCLK_posedge(3),
          TestSignal => PLLCE_PLLCLK_dly(3),
          TestSignalName => "PLLCE(1)",
          TestDelay => tisd_PLLCE_PLLCLK(3),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_PLLCE_PLLCLK_posedge_posedge(3),
          HoldHigh => thold_PLLCE_PLLCLK_posedge_posedge(3),
          SetupLow => tsetup_PLLCE_PLLCLK_negedge_posedge(3),
          HoldLow => thold_PLLCE_PLLCLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_PLLLOCK_PLLCLK_posedge(0),
          TimingData => Tmkr_PLLLOCK_PLLCLK_posedge(0),
          TestSignal => PLLLOCK_PLLCLK_dly(0),
          TestSignalName => "PLLLOCK",
          TestDelay => tisd_PLLLOCK_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_PLLLOCK_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_PLLLOCK_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_PLLLOCK_PLLCLK_negedge_posedge(0),
          HoldLow => thold_PLLLOCK_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
       VitalSetupHoldCheck
        (
          Violation => Tviol_PLLLOCK_PLLCLK_posedge(1),
          TimingData => Tmkr_PLLLOCK_PLLCLK_posedge(1),
          TestSignal => PLLLOCK_PLLCLK_dly(1),
          TestSignalName => "PLLLOCK",
          TestDelay => tisd_PLLLOCK_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_PLLLOCK_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_PLLLOCK_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_PLLLOCK_PLLCLK_negedge_posedge(1),
          HoldLow => thold_PLLLOCK_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
       VitalSetupHoldCheck
        (
          Violation => Tviol_RECAL_PLLCLK_posedge(0),
          TimingData => Tmkr_RECAL_PLLCLK_posedge(0),
          TestSignal => RECAL_PLLCLK_dly(0),
          TestSignalName => "RECAL",
          TestDelay => tisd_RECAL_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_RECAL_PLLCLK_posedge_posedge(0),
          HoldHigh => thold_RECAL_PLLCLK_posedge_posedge(0),
          SetupLow => tsetup_RECAL_PLLCLK_negedge_posedge(0),
          HoldLow => thold_RECAL_PLLCLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_RECAL_PLLCLK_posedge(1),
          TimingData => Tmkr_RECAL_PLLCLK_posedge(1),
          TestSignal => RECAL_PLLCLK_dly(1),
          TestSignalName => "RECAL",
          TestDelay => tisd_RECAL_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_RECAL_PLLCLK_posedge_posedge(1),
          HoldHigh => thold_RECAL_PLLCLK_posedge_posedge(1),
          SetupLow => tsetup_RECAL_PLLCLK_negedge_posedge(1),
          HoldLow => thold_RECAL_PLLCLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_SELFREFRESHENTER_PLLCLK_negedge(0),
          TimingData => Tmkr_SELFREFRESHENTER_PLLCLK_negedge(0),
          TestSignal => SELFREFRESHENTER_PLLCLK_dly(0),
          TestSignalName => "SELFREFRESHENTER",
          TestDelay => tisd_SELFREFRESHENTER_PLLCLK(0),
          RefSignal => PLLCLK_0,
          RefSignalName => "PLLCLK_0",
          RefDelay => ticd_PLLCLK(0),
          SetupHigh => tsetup_SELFREFRESHENTER_PLLCLK_posedge_negedge(0),
          HoldHigh => thold_SELFREFRESHENTER_PLLCLK_posedge_negedge(0),
          SetupLow => tsetup_SELFREFRESHENTER_PLLCLK_negedge_negedge(0),
          HoldLow => thold_SELFREFRESHENTER_PLLCLK_negedge_negedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
         VitalSetupHoldCheck
        (
          Violation => Tviol_SELFREFRESHENTER_PLLCLK_negedge(1),
          TimingData => Tmkr_SELFREFRESHENTER_PLLCLK_negedge(1),
          TestSignal => SELFREFRESHENTER_PLLCLK_dly(1),
          TestSignalName => "SELFREFRESHENTER",
          TestDelay => tisd_SELFREFRESHENTER_PLLCLK(1),
          RefSignal => PLLCLK_1,
          RefSignalName => "PLLCLK_1",
          RefDelay => ticd_PLLCLK(1),
          SetupHigh => tsetup_SELFREFRESHENTER_PLLCLK_posedge_negedge(1),
          HoldHigh => thold_SELFREFRESHENTER_PLLCLK_posedge_negedge(1),
          SetupLow => tsetup_SELFREFRESHENTER_PLLCLK_negedge_negedge(1),
          HoldLow => thold_SELFREFRESHENTER_PLLCLK_negedge_negedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIADDR_UICLK_posedge(0),
          TimingData => Tmkr_UIADDR_UICLK_posedge(0),
          TestSignal => UIADDR_UICLK_dly(0),
          TestSignalName => "UIADDR(0)",
          TestDelay => tisd_UIADDR_UICLK(0),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIADDR_UICLK_posedge_posedge(0),
          HoldHigh => thold_UIADDR_UICLK_posedge_posedge(0),
          SetupLow => tsetup_UIADDR_UICLK_negedge_posedge(0),
          HoldLow => thold_UIADDR_UICLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIADDR_UICLK_posedge(1),
          TimingData => Tmkr_UIADDR_UICLK_posedge(1),
          TestSignal => UIADDR_UICLK_dly(1),
          TestSignalName => "UIADDR(1)",
          TestDelay => tisd_UIADDR_UICLK(1),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIADDR_UICLK_posedge_posedge(1),
          HoldHigh => thold_UIADDR_UICLK_posedge_posedge(1),
          SetupLow => tsetup_UIADDR_UICLK_negedge_posedge(1),
          HoldLow => thold_UIADDR_UICLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIADDR_UICLK_posedge(2),
          TimingData => Tmkr_UIADDR_UICLK_posedge(2),
          TestSignal => UIADDR_UICLK_dly(2),
          TestSignalName => "UIADDR(2)",
          TestDelay => tisd_UIADDR_UICLK(2),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIADDR_UICLK_posedge_posedge(2),
          HoldHigh => thold_UIADDR_UICLK_posedge_posedge(2),
          SetupLow => tsetup_UIADDR_UICLK_negedge_posedge(2),
          HoldLow => thold_UIADDR_UICLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIADDR_UICLK_posedge(3),
          TimingData => Tmkr_UIADDR_UICLK_posedge(3),
          TestSignal => UIADDR_UICLK_dly(3),
          TestSignalName => "UIADDR(3)",
          TestDelay => tisd_UIADDR_UICLK(3),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIADDR_UICLK_posedge_posedge(3),
          HoldHigh => thold_UIADDR_UICLK_posedge_posedge(3),
          SetupLow => tsetup_UIADDR_UICLK_negedge_posedge(3),
          HoldLow => thold_UIADDR_UICLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIADDR_UICLK_posedge(4),
          TimingData => Tmkr_UIADDR_UICLK_posedge(4),
          TestSignal => UIADDR_UICLK_dly(4),
          TestSignalName => "UIADDR(4)",
          TestDelay => tisd_UIADDR_UICLK(4),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIADDR_UICLK_posedge_posedge(4),
          HoldHigh => thold_UIADDR_UICLK_posedge_posedge(4),
          SetupLow => tsetup_UIADDR_UICLK_negedge_posedge(4),
          HoldLow => thold_UIADDR_UICLK_negedge_posedge(4),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIADD_UICLK_posedge,
          TimingData => Tmkr_UIADD_UICLK_posedge,
          TestSignal => UIADD_UICLK_dly,
          TestSignalName => "UIADD",
          TestDelay => tisd_UIADD_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIADD_UICLK_posedge_posedge,
          HoldHigh => thold_UIADD_UICLK_posedge_posedge,
          SetupLow => tsetup_UIADD_UICLK_negedge_posedge,
          HoldLow => thold_UIADD_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIBROADCAST_UICLK_posedge,
          TimingData => Tmkr_UIBROADCAST_UICLK_posedge,
          TestSignal => UIBROADCAST_UICLK_dly,
          TestSignalName => "UIBROADCAST",
          TestDelay => tisd_UIBROADCAST_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIBROADCAST_UICLK_posedge_posedge,
          HoldHigh => thold_UIBROADCAST_UICLK_posedge_posedge,
          SetupLow => tsetup_UIBROADCAST_UICLK_negedge_posedge,
          HoldLow => thold_UIBROADCAST_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UICMDEN_UICLK_posedge,
          TimingData => Tmkr_UICMDEN_UICLK_posedge,
          TestSignal => UICMDEN_UICLK_dly,
          TestSignalName => "UICMDEN",
          TestDelay => tisd_UICMDEN_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UICMDEN_UICLK_posedge_posedge,
          HoldHigh => thold_UICMDEN_UICLK_posedge_posedge,
          SetupLow => tsetup_UICMDEN_UICLK_negedge_posedge,
          HoldLow => thold_UICMDEN_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UICMDIN_UICLK_posedge,
          TimingData => Tmkr_UICMDIN_UICLK_posedge,
          TestSignal => UICMDIN_UICLK_dly,
          TestSignalName => "UICMDIN",
          TestDelay => tisd_UICMDIN_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UICMDIN_UICLK_posedge_posedge,
          HoldHigh => thold_UICMDIN_UICLK_posedge_posedge,
          SetupLow => tsetup_UICMDIN_UICLK_negedge_posedge,
          HoldLow => thold_UICMDIN_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UICMD_UICLK_posedge,
          TimingData => Tmkr_UICMD_UICLK_posedge,
          TestSignal => UICMD_UICLK_dly,
          TestSignalName => "UICMD",
          TestDelay => tisd_UICMD_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UICMD_UICLK_posedge_posedge,
          HoldHigh => thold_UICMD_UICLK_posedge_posedge,
          SetupLow => tsetup_UICMD_UICLK_negedge_posedge,
          HoldLow => thold_UICMD_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UICS_UICLK_posedge,
          TimingData => Tmkr_UICS_UICLK_posedge,
          TestSignal => UICS_UICLK_dly,
          TestSignalName => "UICS",
          TestDelay => tisd_UICS_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UICS_UICLK_posedge_posedge,
          HoldHigh => thold_UICS_UICLK_posedge_posedge,
          SetupLow => tsetup_UICS_UICLK_negedge_posedge,
          HoldLow => thold_UICS_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDONECAL_UICLK_posedge,
          TimingData => Tmkr_UIDONECAL_UICLK_posedge,
          TestSignal => UIDONECAL_UICLK_dly,
          TestSignalName => "UIDONECAL",
          TestDelay => tisd_UIDONECAL_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDONECAL_UICLK_posedge_posedge,
          HoldHigh => thold_UIDONECAL_UICLK_posedge_posedge,
          SetupLow => tsetup_UIDONECAL_UICLK_negedge_posedge,
          HoldLow => thold_UIDONECAL_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQCOUNT_UICLK_posedge(0),
          TimingData => Tmkr_UIDQCOUNT_UICLK_posedge(0),
          TestSignal => UIDQCOUNT_UICLK_dly(0),
          TestSignalName => "UIDQCOUNT(0)",
          TestDelay => tisd_UIDQCOUNT_UICLK(0),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQCOUNT_UICLK_posedge_posedge(0),
          HoldHigh => thold_UIDQCOUNT_UICLK_posedge_posedge(0),
          SetupLow => tsetup_UIDQCOUNT_UICLK_negedge_posedge(0),
          HoldLow => thold_UIDQCOUNT_UICLK_negedge_posedge(0),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQCOUNT_UICLK_posedge(1),
          TimingData => Tmkr_UIDQCOUNT_UICLK_posedge(1),
          TestSignal => UIDQCOUNT_UICLK_dly(1),
          TestSignalName => "UIDQCOUNT(1)",
          TestDelay => tisd_UIDQCOUNT_UICLK(1),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQCOUNT_UICLK_posedge_posedge(1),
          HoldHigh => thold_UIDQCOUNT_UICLK_posedge_posedge(1),
          SetupLow => tsetup_UIDQCOUNT_UICLK_negedge_posedge(1),
          HoldLow => thold_UIDQCOUNT_UICLK_negedge_posedge(1),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQCOUNT_UICLK_posedge(2),
          TimingData => Tmkr_UIDQCOUNT_UICLK_posedge(2),
          TestSignal => UIDQCOUNT_UICLK_dly(2),
          TestSignalName => "UIDQCOUNT(2)",
          TestDelay => tisd_UIDQCOUNT_UICLK(2),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQCOUNT_UICLK_posedge_posedge(2),
          HoldHigh => thold_UIDQCOUNT_UICLK_posedge_posedge(2),
          SetupLow => tsetup_UIDQCOUNT_UICLK_negedge_posedge(2),
          HoldLow => thold_UIDQCOUNT_UICLK_negedge_posedge(2),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQCOUNT_UICLK_posedge(3),
          TimingData => Tmkr_UIDQCOUNT_UICLK_posedge(3),
          TestSignal => UIDQCOUNT_UICLK_dly(3),
          TestSignalName => "UIDQCOUNT(3)",
          TestDelay => tisd_UIDQCOUNT_UICLK(3),
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQCOUNT_UICLK_posedge_posedge(3),
          HoldHigh => thold_UIDQCOUNT_UICLK_posedge_posedge(3),
          SetupLow => tsetup_UIDQCOUNT_UICLK_negedge_posedge(3),
          HoldLow => thold_UIDQCOUNT_UICLK_negedge_posedge(3),
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQLOWERDEC_UICLK_posedge,
          TimingData => Tmkr_UIDQLOWERDEC_UICLK_posedge,
          TestSignal => UIDQLOWERDEC_UICLK_dly,
          TestSignalName => "UIDQLOWERDEC",
          TestDelay => tisd_UIDQLOWERDEC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQLOWERDEC_UICLK_posedge_posedge,
          HoldHigh => thold_UIDQLOWERDEC_UICLK_posedge_posedge,
          SetupLow => tsetup_UIDQLOWERDEC_UICLK_negedge_posedge,
          HoldLow => thold_UIDQLOWERDEC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQLOWERINC_UICLK_posedge,
          TimingData => Tmkr_UIDQLOWERINC_UICLK_posedge,
          TestSignal => UIDQLOWERINC_UICLK_dly,
          TestSignalName => "UIDQLOWERINC",
          TestDelay => tisd_UIDQLOWERINC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQLOWERINC_UICLK_posedge_posedge,
          HoldHigh => thold_UIDQLOWERINC_UICLK_posedge_posedge,
          SetupLow => tsetup_UIDQLOWERINC_UICLK_negedge_posedge,
          HoldLow => thold_UIDQLOWERINC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQUPPERDEC_UICLK_posedge,
          TimingData => Tmkr_UIDQUPPERDEC_UICLK_posedge,
          TestSignal => UIDQUPPERDEC_UICLK_dly,
          TestSignalName => "UIDQUPPERDEC",
          TestDelay => tisd_UIDQUPPERDEC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQUPPERDEC_UICLK_posedge_posedge,
          HoldHigh => thold_UIDQUPPERDEC_UICLK_posedge_posedge,
          SetupLow => tsetup_UIDQUPPERDEC_UICLK_negedge_posedge,
          HoldLow => thold_UIDQUPPERDEC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDQUPPERINC_UICLK_posedge,
          TimingData => Tmkr_UIDQUPPERINC_UICLK_posedge,
          TestSignal => UIDQUPPERINC_UICLK_dly,
          TestSignalName => "UIDQUPPERINC",
          TestDelay => tisd_UIDQUPPERINC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDQUPPERINC_UICLK_posedge_posedge,
          HoldHigh => thold_UIDQUPPERINC_UICLK_posedge_posedge,
          SetupLow => tsetup_UIDQUPPERINC_UICLK_negedge_posedge,
          HoldLow => thold_UIDQUPPERINC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIDRPUPDATE_UICLK_posedge,
          TimingData => Tmkr_UIDRPUPDATE_UICLK_posedge,
          TestSignal => UIDRPUPDATE_UICLK_dly,
          TestSignalName => "UIDRPUPDATE",
          TestDelay => tisd_UIDRPUPDATE_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIDRPUPDATE_UICLK_posedge_posedge,
          HoldHigh => thold_UIDRPUPDATE_UICLK_posedge_posedge,
          SetupLow => tsetup_UIDRPUPDATE_UICLK_negedge_posedge,
          HoldLow => thold_UIDRPUPDATE_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UILDQSDEC_UICLK_posedge,
          TimingData => Tmkr_UILDQSDEC_UICLK_posedge,
          TestSignal => UILDQSDEC_UICLK_dly,
          TestSignalName => "UILDQSDEC",
          TestDelay => tisd_UILDQSDEC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UILDQSDEC_UICLK_posedge_posedge,
          HoldHigh => thold_UILDQSDEC_UICLK_posedge_posedge,
          SetupLow => tsetup_UILDQSDEC_UICLK_negedge_posedge,
          HoldLow => thold_UILDQSDEC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UILDQSINC_UICLK_posedge,
          TimingData => Tmkr_UILDQSINC_UICLK_posedge,
          TestSignal => UILDQSINC_UICLK_dly,
          TestSignalName => "UILDQSINC",
          TestDelay => tisd_UILDQSINC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UILDQSINC_UICLK_posedge_posedge,
          HoldHigh => thold_UILDQSINC_UICLK_posedge_posedge,
          SetupLow => tsetup_UILDQSINC_UICLK_negedge_posedge,
          HoldLow => thold_UILDQSINC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIREAD_UICLK_posedge,
          TimingData => Tmkr_UIREAD_UICLK_posedge,
          TestSignal => UIREAD_UICLK_dly,
          TestSignalName => "UIREAD",
          TestDelay => tisd_UIREAD_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIREAD_UICLK_posedge_posedge,
          HoldHigh => thold_UIREAD_UICLK_posedge_posedge,
          SetupLow => tsetup_UIREAD_UICLK_negedge_posedge,
          HoldLow => thold_UIREAD_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UISDI_UICLK_posedge,
          TimingData => Tmkr_UISDI_UICLK_posedge,
          TestSignal => UISDI_UICLK_dly,
          TestSignalName => "UISDI",
          TestDelay => tisd_UISDI_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UISDI_UICLK_posedge_posedge,
          HoldHigh => thold_UISDI_UICLK_posedge_posedge,
          SetupLow => tsetup_UISDI_UICLK_negedge_posedge,
          HoldLow => thold_UISDI_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIUDQSDEC_UICLK_posedge,
          TimingData => Tmkr_UIUDQSDEC_UICLK_posedge,
          TestSignal => UIUDQSDEC_UICLK_dly,
          TestSignalName => "UIUDQSDEC",
          TestDelay => tisd_UIUDQSDEC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIUDQSDEC_UICLK_posedge_posedge,
          HoldHigh => thold_UIUDQSDEC_UICLK_posedge_posedge,
          SetupLow => tsetup_UIUDQSDEC_UICLK_negedge_posedge,
          HoldLow => thold_UIUDQSDEC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalSetupHoldCheck
        (
          Violation => Tviol_UIUDQSINC_UICLK_posedge,
          TimingData => Tmkr_UIUDQSINC_UICLK_posedge,
          TestSignal => UIUDQSINC_UICLK_dly,
          TestSignalName => "UIUDQSINC",
          TestDelay => tisd_UIUDQSINC_UICLK,
          RefSignal => UICLK_dly,
          RefSignalName => "UICLK",
          RefDelay => ticd_UICLK,
          SetupHigh => tsetup_UIUDQSINC_UICLK_posedge_posedge,
          HoldHigh => thold_UIUDQSINC_UICLK_posedge_posedge,
          SetupLow => tsetup_UIUDQSINC_UICLK_negedge_posedge,
          HoldLow => thold_UIUDQSINC_UICLK_negedge_posedge,
          CheckEnabled   => TRUE,
          RefTransition  => 'R',
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
      end if;
       VitalPathDelay01
        (
          OutSignal     => DQIOWEN0,
          GlitchData    => DQIOWEN0_GlitchData,
          OutSignalName => "DQIOWEN0",
          OutTemp       => DQIOWEN0_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_DQIOWEN0(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );

        VitalPathDelay01
        (
          OutSignal     => DQIOWEN0,
          GlitchData    => DQIOWEN0_GlitchData,
          OutSignalName => "DQIOWEN0",
          OutTemp       => DQIOWEN0_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_DQIOWEN0(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => DQSIOWEN90N,
          GlitchData    => DQSIOWEN90N_GlitchData,
          OutSignalName => "DQSIOWEN90N",
          OutTemp       => DQSIOWEN90N_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_DQSIOWEN90N(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
       VitalPathDelay01
        (
          OutSignal     => DQSIOWEN90N,
          GlitchData    => DQSIOWEN90N_GlitchData,
          OutSignalName => "DQSIOWEN90N",
          OutTemp       => DQSIOWEN90N_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_DQSIOWEN90N(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => DQSIOWEN90P,
          GlitchData    => DQSIOWEN90P_GlitchData,
          OutSignalName => "DQSIOWEN90P",
          OutTemp       => DQSIOWEN90P_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_DQSIOWEN90P(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => DQSIOWEN90P,
          GlitchData    => DQSIOWEN90P_GlitchData,
          OutSignalName => "DQSIOWEN90P",
          OutTemp       => DQSIOWEN90P_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_DQSIOWEN90P(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPADD,
          GlitchData    => IOIDRPADD_GlitchData,
          OutSignalName => "IOIDRPADD",
          OutTemp       => IOIDRPADD_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPADD,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPADDR(0),
          GlitchData    => IOIDRPADDR0_GlitchData,
          OutSignalName => "IOIDRPADDR(0)",
          OutTemp       => IOIDRPADDR_out(0),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPADDR(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPADDR(1),
          GlitchData    => IOIDRPADDR1_GlitchData,
          OutSignalName => "IOIDRPADDR(1)",
          OutTemp       => IOIDRPADDR_out(1),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPADDR(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPADDR(2),
          GlitchData    => IOIDRPADDR2_GlitchData,
          OutSignalName => "IOIDRPADDR(2)",
          OutTemp       => IOIDRPADDR_out(2),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPADDR(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPADDR(3),
          GlitchData    => IOIDRPADDR3_GlitchData,
          OutSignalName => "IOIDRPADDR(3)",
          OutTemp       => IOIDRPADDR_out(3),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPADDR(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPADDR(4),
          GlitchData    => IOIDRPADDR4_GlitchData,
          OutSignalName => "IOIDRPADDR(4)",
          OutTemp       => IOIDRPADDR_out(4),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPADDR(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPBROADCAST,
          GlitchData    => IOIDRPBROADCAST_GlitchData,
          OutSignalName => "IOIDRPBROADCAST",
          OutTemp       => IOIDRPBROADCAST_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPBROADCAST,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPCLK,
          GlitchData    => IOIDRPCLK_GlitchData,
          OutSignalName => "IOIDRPCLK",
          OutTemp       => IOIDRPCLK_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPCLK,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPCS,
          GlitchData    => IOIDRPCS_GlitchData,
          OutSignalName => "IOIDRPCS",
          OutTemp       => IOIDRPCS_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPCS,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPSDO,
          GlitchData    => IOIDRPSDO_GlitchData,
          OutSignalName => "IOIDRPSDO",
          OutTemp       => IOIDRPSDO_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPSDO,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => IOIDRPUPDATE,
          GlitchData    => IOIDRPUPDATE_GlitchData,
          OutSignalName => "IOIDRPUPDATE",
          OutTemp       => IOIDRPUPDATE_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_IOIDRPUPDATE,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0CMDEMPTY,
          GlitchData    => P0CMDEMPTY_GlitchData,
          OutSignalName => "P0CMDEMPTY",
          OutTemp       => P0CMDEMPTY_out,
          Paths       => (0 => (P0CMDCLK_dly'last_event, tpd_P0CMDCLK_P0CMDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0CMDFULL,
          GlitchData    => P0CMDFULL_GlitchData,
          OutSignalName => "P0CMDFULL",
          OutTemp       => P0CMDFULL_out,
          Paths       => (0 => (P0CMDCLK_dly'last_event, tpd_P0CMDCLK_P0CMDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(0),
          GlitchData    => P0RDCOUNT0_GlitchData,
          OutSignalName => "P0RDCOUNT(0)",
          OutTemp       => P0RDCOUNT_out(0),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(1),
          GlitchData    => P0RDCOUNT1_GlitchData,
          OutSignalName => "P0RDCOUNT(1)",
          OutTemp       => P0RDCOUNT_out(1),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(2),
          GlitchData    => P0RDCOUNT2_GlitchData,
          OutSignalName => "P0RDCOUNT(2)",
          OutTemp       => P0RDCOUNT_out(2),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(3),
          GlitchData    => P0RDCOUNT3_GlitchData,
          OutSignalName => "P0RDCOUNT(3)",
          OutTemp       => P0RDCOUNT_out(3),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(4),
          GlitchData    => P0RDCOUNT4_GlitchData,
          OutSignalName => "P0RDCOUNT(4)",
          OutTemp       => P0RDCOUNT_out(4),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(5),
          GlitchData    => P0RDCOUNT5_GlitchData,
          OutSignalName => "P0RDCOUNT(5)",
          OutTemp       => P0RDCOUNT_out(5),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDCOUNT(6),
          GlitchData    => P0RDCOUNT6_GlitchData,
          OutSignalName => "P0RDCOUNT(6)",
          OutTemp       => P0RDCOUNT_out(6),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDCOUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(0),
          GlitchData    => P0RDDATA0_GlitchData,
          OutSignalName => "P0RDDATA(0)",
          OutTemp       => P0RDDATA_out(0),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(1),
          GlitchData    => P0RDDATA1_GlitchData,
          OutSignalName => "P0RDDATA(1)",
          OutTemp       => P0RDDATA_out(1),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(10),
          GlitchData    => P0RDDATA10_GlitchData,
          OutSignalName => "P0RDDATA(10)",
          OutTemp       => P0RDDATA_out(10),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(10),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(11),
          GlitchData    => P0RDDATA11_GlitchData,
          OutSignalName => "P0RDDATA(11)",
          OutTemp       => P0RDDATA_out(11),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(11),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(12),
          GlitchData    => P0RDDATA12_GlitchData,
          OutSignalName => "P0RDDATA(12)",
          OutTemp       => P0RDDATA_out(12),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(12),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(13),
          GlitchData    => P0RDDATA13_GlitchData,
          OutSignalName => "P0RDDATA(13)",
          OutTemp       => P0RDDATA_out(13),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(13),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(14),
          GlitchData    => P0RDDATA14_GlitchData,
          OutSignalName => "P0RDDATA(14)",
          OutTemp       => P0RDDATA_out(14),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(14),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(15),
          GlitchData    => P0RDDATA15_GlitchData,
          OutSignalName => "P0RDDATA(15)",
          OutTemp       => P0RDDATA_out(15),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(15),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(16),
          GlitchData    => P0RDDATA16_GlitchData,
          OutSignalName => "P0RDDATA(16)",
          OutTemp       => P0RDDATA_out(16),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(16),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(17),
          GlitchData    => P0RDDATA17_GlitchData,
          OutSignalName => "P0RDDATA(17)",
          OutTemp       => P0RDDATA_out(17),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(17),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(18),
          GlitchData    => P0RDDATA18_GlitchData,
          OutSignalName => "P0RDDATA(18)",
          OutTemp       => P0RDDATA_out(18),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(18),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(19),
          GlitchData    => P0RDDATA19_GlitchData,
          OutSignalName => "P0RDDATA(19)",
          OutTemp       => P0RDDATA_out(19),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(19),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(2),
          GlitchData    => P0RDDATA2_GlitchData,
          OutSignalName => "P0RDDATA(2)",
          OutTemp       => P0RDDATA_out(2),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(20),
          GlitchData    => P0RDDATA20_GlitchData,
          OutSignalName => "P0RDDATA(20)",
          OutTemp       => P0RDDATA_out(20),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(20),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(21),
          GlitchData    => P0RDDATA21_GlitchData,
          OutSignalName => "P0RDDATA(21)",
          OutTemp       => P0RDDATA_out(21),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(21),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(22),
          GlitchData    => P0RDDATA22_GlitchData,
          OutSignalName => "P0RDDATA(22)",
          OutTemp       => P0RDDATA_out(22),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(22),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(23),
          GlitchData    => P0RDDATA23_GlitchData,
          OutSignalName => "P0RDDATA(23)",
          OutTemp       => P0RDDATA_out(23),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(23),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(24),
          GlitchData    => P0RDDATA24_GlitchData,
          OutSignalName => "P0RDDATA(24)",
          OutTemp       => P0RDDATA_out(24),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(24),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(25),
          GlitchData    => P0RDDATA25_GlitchData,
          OutSignalName => "P0RDDATA(25)",
          OutTemp       => P0RDDATA_out(25),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(25),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(26),
          GlitchData    => P0RDDATA26_GlitchData,
          OutSignalName => "P0RDDATA(26)",
          OutTemp       => P0RDDATA_out(26),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(26),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(27),
          GlitchData    => P0RDDATA27_GlitchData,
          OutSignalName => "P0RDDATA(27)",
          OutTemp       => P0RDDATA_out(27),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(27),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(28),
          GlitchData    => P0RDDATA28_GlitchData,
          OutSignalName => "P0RDDATA(28)",
          OutTemp       => P0RDDATA_out(28),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(28),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(29),
          GlitchData    => P0RDDATA29_GlitchData,
          OutSignalName => "P0RDDATA(29)",
          OutTemp       => P0RDDATA_out(29),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(29),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(3),
          GlitchData    => P0RDDATA3_GlitchData,
          OutSignalName => "P0RDDATA(3)",
          OutTemp       => P0RDDATA_out(3),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(30),
          GlitchData    => P0RDDATA30_GlitchData,
          OutSignalName => "P0RDDATA(30)",
          OutTemp       => P0RDDATA_out(30),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(30),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(31),
          GlitchData    => P0RDDATA31_GlitchData,
          OutSignalName => "P0RDDATA(31)",
          OutTemp       => P0RDDATA_out(31),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(31),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(4),
          GlitchData    => P0RDDATA4_GlitchData,
          OutSignalName => "P0RDDATA(4)",
          OutTemp       => P0RDDATA_out(4),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(5),
          GlitchData    => P0RDDATA5_GlitchData,
          OutSignalName => "P0RDDATA(5)",
          OutTemp       => P0RDDATA_out(5),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(6),
          GlitchData    => P0RDDATA6_GlitchData,
          OutSignalName => "P0RDDATA(6)",
          OutTemp       => P0RDDATA_out(6),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(7),
          GlitchData    => P0RDDATA7_GlitchData,
          OutSignalName => "P0RDDATA(7)",
          OutTemp       => P0RDDATA_out(7),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(8),
          GlitchData    => P0RDDATA8_GlitchData,
          OutSignalName => "P0RDDATA(8)",
          OutTemp       => P0RDDATA_out(8),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(8),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDDATA(9),
          GlitchData    => P0RDDATA9_GlitchData,
          OutSignalName => "P0RDDATA(9)",
          OutTemp       => P0RDDATA_out(9),
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDDATA(9),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDEMPTY,
          GlitchData    => P0RDEMPTY_GlitchData,
          OutSignalName => "P0RDEMPTY",
          OutTemp       => P0RDEMPTY_out,
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDERROR,
          GlitchData    => P0RDERROR_GlitchData,
          OutSignalName => "P0RDERROR",
          OutTemp       => P0RDERROR_out,
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDFULL,
          GlitchData    => P0RDFULL_GlitchData,
          OutSignalName => "P0RDFULL",
          OutTemp       => P0RDFULL_out,
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0RDOVERFLOW,
          GlitchData    => P0RDOVERFLOW_GlitchData,
          OutSignalName => "P0RDOVERFLOW",
          OutTemp       => P0RDOVERFLOW_out,
          Paths       => (0 => (P0RDCLK_dly'last_event, tpd_P0RDCLK_P0RDOVERFLOW,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(0),
          GlitchData    => P0WRCOUNT0_GlitchData,
          OutSignalName => "P0WRCOUNT(0)",
          OutTemp       => P0WRCOUNT_out(0),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(1),
          GlitchData    => P0WRCOUNT1_GlitchData,
          OutSignalName => "P0WRCOUNT(1)",
          OutTemp       => P0WRCOUNT_out(1),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(2),
          GlitchData    => P0WRCOUNT2_GlitchData,
          OutSignalName => "P0WRCOUNT(2)",
          OutTemp       => P0WRCOUNT_out(2),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(3),
          GlitchData    => P0WRCOUNT3_GlitchData,
          OutSignalName => "P0WRCOUNT(3)",
          OutTemp       => P0WRCOUNT_out(3),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(4),
          GlitchData    => P0WRCOUNT4_GlitchData,
          OutSignalName => "P0WRCOUNT(4)",
          OutTemp       => P0WRCOUNT_out(4),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(5),
          GlitchData    => P0WRCOUNT5_GlitchData,
          OutSignalName => "P0WRCOUNT(5)",
          OutTemp       => P0WRCOUNT_out(5),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRCOUNT(6),
          GlitchData    => P0WRCOUNT6_GlitchData,
          OutSignalName => "P0WRCOUNT(6)",
          OutTemp       => P0WRCOUNT_out(6),
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRCOUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WREMPTY,
          GlitchData    => P0WREMPTY_GlitchData,
          OutSignalName => "P0WREMPTY",
          OutTemp       => P0WREMPTY_out,
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WREMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRERROR,
          GlitchData    => P0WRERROR_GlitchData,
          OutSignalName => "P0WRERROR",
          OutTemp       => P0WRERROR_out,
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRFULL,
          GlitchData    => P0WRFULL_GlitchData,
          OutSignalName => "P0WRFULL",
          OutTemp       => P0WRFULL_out,
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P0WRUNDERRUN,
          GlitchData    => P0WRUNDERRUN_GlitchData,
          OutSignalName => "P0WRUNDERRUN",
          OutTemp       => P0WRUNDERRUN_out,
          Paths       => (0 => (P0WRCLK_dly'last_event, tpd_P0WRCLK_P0WRUNDERRUN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1CMDEMPTY,
          GlitchData    => P1CMDEMPTY_GlitchData,
          OutSignalName => "P1CMDEMPTY",
          OutTemp       => P1CMDEMPTY_out,
          Paths       => (0 => (P1CMDCLK_dly'last_event, tpd_P1CMDCLK_P1CMDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1CMDFULL,
          GlitchData    => P1CMDFULL_GlitchData,
          OutSignalName => "P1CMDFULL",
          OutTemp       => P1CMDFULL_out,
          Paths       => (0 => (P1CMDCLK_dly'last_event, tpd_P1CMDCLK_P1CMDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(0),
          GlitchData    => P1RDCOUNT0_GlitchData,
          OutSignalName => "P1RDCOUNT(0)",
          OutTemp       => P1RDCOUNT_out(0),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(1),
          GlitchData    => P1RDCOUNT1_GlitchData,
          OutSignalName => "P1RDCOUNT(1)",
          OutTemp       => P1RDCOUNT_out(1),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(2),
          GlitchData    => P1RDCOUNT2_GlitchData,
          OutSignalName => "P1RDCOUNT(2)",
          OutTemp       => P1RDCOUNT_out(2),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(3),
          GlitchData    => P1RDCOUNT3_GlitchData,
          OutSignalName => "P1RDCOUNT(3)",
          OutTemp       => P1RDCOUNT_out(3),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(4),
          GlitchData    => P1RDCOUNT4_GlitchData,
          OutSignalName => "P1RDCOUNT(4)",
          OutTemp       => P1RDCOUNT_out(4),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(5),
          GlitchData    => P1RDCOUNT5_GlitchData,
          OutSignalName => "P1RDCOUNT(5)",
          OutTemp       => P1RDCOUNT_out(5),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDCOUNT(6),
          GlitchData    => P1RDCOUNT6_GlitchData,
          OutSignalName => "P1RDCOUNT(6)",
          OutTemp       => P1RDCOUNT_out(6),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDCOUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(0),
          GlitchData    => P1RDDATA0_GlitchData,
          OutSignalName => "P1RDDATA(0)",
          OutTemp       => P1RDDATA_out(0),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(1),
          GlitchData    => P1RDDATA1_GlitchData,
          OutSignalName => "P1RDDATA(1)",
          OutTemp       => P1RDDATA_out(1),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(10),
          GlitchData    => P1RDDATA10_GlitchData,
          OutSignalName => "P1RDDATA(10)",
          OutTemp       => P1RDDATA_out(10),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(10),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(11),
          GlitchData    => P1RDDATA11_GlitchData,
          OutSignalName => "P1RDDATA(11)",
          OutTemp       => P1RDDATA_out(11),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(11),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(12),
          GlitchData    => P1RDDATA12_GlitchData,
          OutSignalName => "P1RDDATA(12)",
          OutTemp       => P1RDDATA_out(12),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(12),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(13),
          GlitchData    => P1RDDATA13_GlitchData,
          OutSignalName => "P1RDDATA(13)",
          OutTemp       => P1RDDATA_out(13),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(13),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(14),
          GlitchData    => P1RDDATA14_GlitchData,
          OutSignalName => "P1RDDATA(14)",
          OutTemp       => P1RDDATA_out(14),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(14),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(15),
          GlitchData    => P1RDDATA15_GlitchData,
          OutSignalName => "P1RDDATA(15)",
          OutTemp       => P1RDDATA_out(15),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(15),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(16),
          GlitchData    => P1RDDATA16_GlitchData,
          OutSignalName => "P1RDDATA(16)",
          OutTemp       => P1RDDATA_out(16),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(16),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(17),
          GlitchData    => P1RDDATA17_GlitchData,
          OutSignalName => "P1RDDATA(17)",
          OutTemp       => P1RDDATA_out(17),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(17),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(18),
          GlitchData    => P1RDDATA18_GlitchData,
          OutSignalName => "P1RDDATA(18)",
          OutTemp       => P1RDDATA_out(18),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(18),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(19),
          GlitchData    => P1RDDATA19_GlitchData,
          OutSignalName => "P1RDDATA(19)",
          OutTemp       => P1RDDATA_out(19),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(19),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(2),
          GlitchData    => P1RDDATA2_GlitchData,
          OutSignalName => "P1RDDATA(2)",
          OutTemp       => P1RDDATA_out(2),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(20),
          GlitchData    => P1RDDATA20_GlitchData,
          OutSignalName => "P1RDDATA(20)",
          OutTemp       => P1RDDATA_out(20),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(20),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(21),
          GlitchData    => P1RDDATA21_GlitchData,
          OutSignalName => "P1RDDATA(21)",
          OutTemp       => P1RDDATA_out(21),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(21),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(22),
          GlitchData    => P1RDDATA22_GlitchData,
          OutSignalName => "P1RDDATA(22)",
          OutTemp       => P1RDDATA_out(22),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(22),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(23),
          GlitchData    => P1RDDATA23_GlitchData,
          OutSignalName => "P1RDDATA(23)",
          OutTemp       => P1RDDATA_out(23),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(23),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(24),
          GlitchData    => P1RDDATA24_GlitchData,
          OutSignalName => "P1RDDATA(24)",
          OutTemp       => P1RDDATA_out(24),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(24),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(25),
          GlitchData    => P1RDDATA25_GlitchData,
          OutSignalName => "P1RDDATA(25)",
          OutTemp       => P1RDDATA_out(25),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(25),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(26),
          GlitchData    => P1RDDATA26_GlitchData,
          OutSignalName => "P1RDDATA(26)",
          OutTemp       => P1RDDATA_out(26),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(26),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(27),
          GlitchData    => P1RDDATA27_GlitchData,
          OutSignalName => "P1RDDATA(27)",
          OutTemp       => P1RDDATA_out(27),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(27),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(28),
          GlitchData    => P1RDDATA28_GlitchData,
          OutSignalName => "P1RDDATA(28)",
          OutTemp       => P1RDDATA_out(28),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(28),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(29),
          GlitchData    => P1RDDATA29_GlitchData,
          OutSignalName => "P1RDDATA(29)",
          OutTemp       => P1RDDATA_out(29),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(29),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(3),
          GlitchData    => P1RDDATA3_GlitchData,
          OutSignalName => "P1RDDATA(3)",
          OutTemp       => P1RDDATA_out(3),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(30),
          GlitchData    => P1RDDATA30_GlitchData,
          OutSignalName => "P1RDDATA(30)",
          OutTemp       => P1RDDATA_out(30),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(30),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(31),
          GlitchData    => P1RDDATA31_GlitchData,
          OutSignalName => "P1RDDATA(31)",
          OutTemp       => P1RDDATA_out(31),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(31),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(4),
          GlitchData    => P1RDDATA4_GlitchData,
          OutSignalName => "P1RDDATA(4)",
          OutTemp       => P1RDDATA_out(4),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(5),
          GlitchData    => P1RDDATA5_GlitchData,
          OutSignalName => "P1RDDATA(5)",
          OutTemp       => P1RDDATA_out(5),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(6),
          GlitchData    => P1RDDATA6_GlitchData,
          OutSignalName => "P1RDDATA(6)",
          OutTemp       => P1RDDATA_out(6),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(7),
          GlitchData    => P1RDDATA7_GlitchData,
          OutSignalName => "P1RDDATA(7)",
          OutTemp       => P1RDDATA_out(7),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(8),
          GlitchData    => P1RDDATA8_GlitchData,
          OutSignalName => "P1RDDATA(8)",
          OutTemp       => P1RDDATA_out(8),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(8),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDDATA(9),
          GlitchData    => P1RDDATA9_GlitchData,
          OutSignalName => "P1RDDATA(9)",
          OutTemp       => P1RDDATA_out(9),
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDDATA(9),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDEMPTY,
          GlitchData    => P1RDEMPTY_GlitchData,
          OutSignalName => "P1RDEMPTY",
          OutTemp       => P1RDEMPTY_out,
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDERROR,
          GlitchData    => P1RDERROR_GlitchData,
          OutSignalName => "P1RDERROR",
          OutTemp       => P1RDERROR_out,
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDFULL,
          GlitchData    => P1RDFULL_GlitchData,
          OutSignalName => "P1RDFULL",
          OutTemp       => P1RDFULL_out,
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1RDOVERFLOW,
          GlitchData    => P1RDOVERFLOW_GlitchData,
          OutSignalName => "P1RDOVERFLOW",
          OutTemp       => P1RDOVERFLOW_out,
          Paths       => (0 => (P1RDCLK_dly'last_event, tpd_P1RDCLK_P1RDOVERFLOW,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(0),
          GlitchData    => P1WRCOUNT0_GlitchData,
          OutSignalName => "P1WRCOUNT(0)",
          OutTemp       => P1WRCOUNT_out(0),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(1),
          GlitchData    => P1WRCOUNT1_GlitchData,
          OutSignalName => "P1WRCOUNT(1)",
          OutTemp       => P1WRCOUNT_out(1),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(2),
          GlitchData    => P1WRCOUNT2_GlitchData,
          OutSignalName => "P1WRCOUNT(2)",
          OutTemp       => P1WRCOUNT_out(2),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(3),
          GlitchData    => P1WRCOUNT3_GlitchData,
          OutSignalName => "P1WRCOUNT(3)",
          OutTemp       => P1WRCOUNT_out(3),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(4),
          GlitchData    => P1WRCOUNT4_GlitchData,
          OutSignalName => "P1WRCOUNT(4)",
          OutTemp       => P1WRCOUNT_out(4),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(5),
          GlitchData    => P1WRCOUNT5_GlitchData,
          OutSignalName => "P1WRCOUNT(5)",
          OutTemp       => P1WRCOUNT_out(5),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRCOUNT(6),
          GlitchData    => P1WRCOUNT6_GlitchData,
          OutSignalName => "P1WRCOUNT(6)",
          OutTemp       => P1WRCOUNT_out(6),
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRCOUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WREMPTY,
          GlitchData    => P1WREMPTY_GlitchData,
          OutSignalName => "P1WREMPTY",
          OutTemp       => P1WREMPTY_out,
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WREMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRERROR,
          GlitchData    => P1WRERROR_GlitchData,
          OutSignalName => "P1WRERROR",
          OutTemp       => P1WRERROR_out,
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRFULL,
          GlitchData    => P1WRFULL_GlitchData,
          OutSignalName => "P1WRFULL",
          OutTemp       => P1WRFULL_out,
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P1WRUNDERRUN,
          GlitchData    => P1WRUNDERRUN_GlitchData,
          OutSignalName => "P1WRUNDERRUN",
          OutTemp       => P1WRUNDERRUN_out,
          Paths       => (0 => (P1WRCLK_dly'last_event, tpd_P1WRCLK_P1WRUNDERRUN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2CMDEMPTY,
          GlitchData    => P2CMDEMPTY_GlitchData,
          OutSignalName => "P2CMDEMPTY",
          OutTemp       => P2CMDEMPTY_out,
          Paths       => (0 => (P2CMDCLK_dly'last_event, tpd_P2CMDCLK_P2CMDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2CMDFULL,
          GlitchData    => P2CMDFULL_GlitchData,
          OutSignalName => "P2CMDFULL",
          OutTemp       => P2CMDFULL_out,
          Paths       => (0 => (P2CMDCLK_dly'last_event, tpd_P2CMDCLK_P2CMDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(0),
          GlitchData    => P2COUNT0_GlitchData,
          OutSignalName => "P2COUNT(0)",
          OutTemp       => P2COUNT_out(0),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(1),
          GlitchData    => P2COUNT1_GlitchData,
          OutSignalName => "P2COUNT(1)",
          OutTemp       => P2COUNT_out(1),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(2),
          GlitchData    => P2COUNT2_GlitchData,
          OutSignalName => "P2COUNT(2)",
          OutTemp       => P2COUNT_out(2),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(3),
          GlitchData    => P2COUNT3_GlitchData,
          OutSignalName => "P2COUNT(3)",
          OutTemp       => P2COUNT_out(3),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(4),
          GlitchData    => P2COUNT4_GlitchData,
          OutSignalName => "P2COUNT(4)",
          OutTemp       => P2COUNT_out(4),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(5),
          GlitchData    => P2COUNT5_GlitchData,
          OutSignalName => "P2COUNT(5)",
          OutTemp       => P2COUNT_out(5),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2COUNT(6),
          GlitchData    => P2COUNT6_GlitchData,
          OutSignalName => "P2COUNT(6)",
          OutTemp       => P2COUNT_out(6),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2COUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2EMPTY,
          GlitchData    => P2EMPTY_GlitchData,
          OutSignalName => "P2EMPTY",
          OutTemp       => P2EMPTY_out,
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2EMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2ERROR,
          GlitchData    => P2ERROR_GlitchData,
          OutSignalName => "P2ERROR",
          OutTemp       => P2ERROR_out,
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2ERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2FULL,
          GlitchData    => P2FULL_GlitchData,
          OutSignalName => "P2FULL",
          OutTemp       => P2FULL_out,
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2FULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(0),
          GlitchData    => P2RDDATA0_GlitchData,
          OutSignalName => "P2RDDATA(0)",
          OutTemp       => P2RDDATA_out(0),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(1),
          GlitchData    => P2RDDATA1_GlitchData,
          OutSignalName => "P2RDDATA(1)",
          OutTemp       => P2RDDATA_out(1),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(10),
          GlitchData    => P2RDDATA10_GlitchData,
          OutSignalName => "P2RDDATA(10)",
          OutTemp       => P2RDDATA_out(10),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(10),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(11),
          GlitchData    => P2RDDATA11_GlitchData,
          OutSignalName => "P2RDDATA(11)",
          OutTemp       => P2RDDATA_out(11),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(11),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(12),
          GlitchData    => P2RDDATA12_GlitchData,
          OutSignalName => "P2RDDATA(12)",
          OutTemp       => P2RDDATA_out(12),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(12),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(13),
          GlitchData    => P2RDDATA13_GlitchData,
          OutSignalName => "P2RDDATA(13)",
          OutTemp       => P2RDDATA_out(13),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(13),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(14),
          GlitchData    => P2RDDATA14_GlitchData,
          OutSignalName => "P2RDDATA(14)",
          OutTemp       => P2RDDATA_out(14),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(14),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(15),
          GlitchData    => P2RDDATA15_GlitchData,
          OutSignalName => "P2RDDATA(15)",
          OutTemp       => P2RDDATA_out(15),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(15),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(16),
          GlitchData    => P2RDDATA16_GlitchData,
          OutSignalName => "P2RDDATA(16)",
          OutTemp       => P2RDDATA_out(16),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(16),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(17),
          GlitchData    => P2RDDATA17_GlitchData,
          OutSignalName => "P2RDDATA(17)",
          OutTemp       => P2RDDATA_out(17),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(17),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(18),
          GlitchData    => P2RDDATA18_GlitchData,
          OutSignalName => "P2RDDATA(18)",
          OutTemp       => P2RDDATA_out(18),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(18),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(19),
          GlitchData    => P2RDDATA19_GlitchData,
          OutSignalName => "P2RDDATA(19)",
          OutTemp       => P2RDDATA_out(19),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(19),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(2),
          GlitchData    => P2RDDATA2_GlitchData,
          OutSignalName => "P2RDDATA(2)",
          OutTemp       => P2RDDATA_out(2),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(20),
          GlitchData    => P2RDDATA20_GlitchData,
          OutSignalName => "P2RDDATA(20)",
          OutTemp       => P2RDDATA_out(20),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(20),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(21),
          GlitchData    => P2RDDATA21_GlitchData,
          OutSignalName => "P2RDDATA(21)",
          OutTemp       => P2RDDATA_out(21),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(21),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(22),
          GlitchData    => P2RDDATA22_GlitchData,
          OutSignalName => "P2RDDATA(22)",
          OutTemp       => P2RDDATA_out(22),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(22),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(23),
          GlitchData    => P2RDDATA23_GlitchData,
          OutSignalName => "P2RDDATA(23)",
          OutTemp       => P2RDDATA_out(23),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(23),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(24),
          GlitchData    => P2RDDATA24_GlitchData,
          OutSignalName => "P2RDDATA(24)",
          OutTemp       => P2RDDATA_out(24),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(24),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(25),
          GlitchData    => P2RDDATA25_GlitchData,
          OutSignalName => "P2RDDATA(25)",
          OutTemp       => P2RDDATA_out(25),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(25),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(26),
          GlitchData    => P2RDDATA26_GlitchData,
          OutSignalName => "P2RDDATA(26)",
          OutTemp       => P2RDDATA_out(26),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(26),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(27),
          GlitchData    => P2RDDATA27_GlitchData,
          OutSignalName => "P2RDDATA(27)",
          OutTemp       => P2RDDATA_out(27),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(27),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(28),
          GlitchData    => P2RDDATA28_GlitchData,
          OutSignalName => "P2RDDATA(28)",
          OutTemp       => P2RDDATA_out(28),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(28),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(29),
          GlitchData    => P2RDDATA29_GlitchData,
          OutSignalName => "P2RDDATA(29)",
          OutTemp       => P2RDDATA_out(29),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(29),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(3),
          GlitchData    => P2RDDATA3_GlitchData,
          OutSignalName => "P2RDDATA(3)",
          OutTemp       => P2RDDATA_out(3),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(30),
          GlitchData    => P2RDDATA30_GlitchData,
          OutSignalName => "P2RDDATA(30)",
          OutTemp       => P2RDDATA_out(30),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(30),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(31),
          GlitchData    => P2RDDATA31_GlitchData,
          OutSignalName => "P2RDDATA(31)",
          OutTemp       => P2RDDATA_out(31),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(31),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(4),
          GlitchData    => P2RDDATA4_GlitchData,
          OutSignalName => "P2RDDATA(4)",
          OutTemp       => P2RDDATA_out(4),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(5),
          GlitchData    => P2RDDATA5_GlitchData,
          OutSignalName => "P2RDDATA(5)",
          OutTemp       => P2RDDATA_out(5),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(6),
          GlitchData    => P2RDDATA6_GlitchData,
          OutSignalName => "P2RDDATA(6)",
          OutTemp       => P2RDDATA_out(6),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(7),
          GlitchData    => P2RDDATA7_GlitchData,
          OutSignalName => "P2RDDATA(7)",
          OutTemp       => P2RDDATA_out(7),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(8),
          GlitchData    => P2RDDATA8_GlitchData,
          OutSignalName => "P2RDDATA(8)",
          OutTemp       => P2RDDATA_out(8),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(8),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDDATA(9),
          GlitchData    => P2RDDATA9_GlitchData,
          OutSignalName => "P2RDDATA(9)",
          OutTemp       => P2RDDATA_out(9),
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDDATA(9),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2RDOVERFLOW,
          GlitchData    => P2RDOVERFLOW_GlitchData,
          OutSignalName => "P2RDOVERFLOW",
          OutTemp       => P2RDOVERFLOW_out,
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2RDOVERFLOW,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P2WRUNDERRUN,
          GlitchData    => P2WRUNDERRUN_GlitchData,
          OutSignalName => "P2WRUNDERRUN",
          OutTemp       => P2WRUNDERRUN_out,
          Paths       => (0 => (P2CLK_dly'last_event, tpd_P2CLK_P2WRUNDERRUN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3CMDEMPTY,
          GlitchData    => P3CMDEMPTY_GlitchData,
          OutSignalName => "P3CMDEMPTY",
          OutTemp       => P3CMDEMPTY_out,
          Paths       => (0 => (P3CMDCLK_dly'last_event, tpd_P3CMDCLK_P3CMDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3CMDFULL,
          GlitchData    => P3CMDFULL_GlitchData,
          OutSignalName => "P3CMDFULL",
          OutTemp       => P3CMDFULL_out,
          Paths       => (0 => (P3CMDCLK_dly'last_event, tpd_P3CMDCLK_P3CMDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(0),
          GlitchData    => P3COUNT0_GlitchData,
          OutSignalName => "P3COUNT(0)",
          OutTemp       => P3COUNT_out(0),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(1),
          GlitchData    => P3COUNT1_GlitchData,
          OutSignalName => "P3COUNT(1)",
          OutTemp       => P3COUNT_out(1),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(2),
          GlitchData    => P3COUNT2_GlitchData,
          OutSignalName => "P3COUNT(2)",
          OutTemp       => P3COUNT_out(2),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(3),
          GlitchData    => P3COUNT3_GlitchData,
          OutSignalName => "P3COUNT(3)",
          OutTemp       => P3COUNT_out(3),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(4),
          GlitchData    => P3COUNT4_GlitchData,
          OutSignalName => "P3COUNT(4)",
          OutTemp       => P3COUNT_out(4),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(5),
          GlitchData    => P3COUNT5_GlitchData,
          OutSignalName => "P3COUNT(5)",
          OutTemp       => P3COUNT_out(5),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3COUNT(6),
          GlitchData    => P3COUNT6_GlitchData,
          OutSignalName => "P3COUNT(6)",
          OutTemp       => P3COUNT_out(6),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3COUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3EMPTY,
          GlitchData    => P3EMPTY_GlitchData,
          OutSignalName => "P3EMPTY",
          OutTemp       => P3EMPTY_out,
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3EMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3ERROR,
          GlitchData    => P3ERROR_GlitchData,
          OutSignalName => "P3ERROR",
          OutTemp       => P3ERROR_out,
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3ERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3FULL,
          GlitchData    => P3FULL_GlitchData,
          OutSignalName => "P3FULL",
          OutTemp       => P3FULL_out,
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3FULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(0),
          GlitchData    => P3RDDATA0_GlitchData,
          OutSignalName => "P3RDDATA(0)",
          OutTemp       => P3RDDATA_out(0),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(1),
          GlitchData    => P3RDDATA1_GlitchData,
          OutSignalName => "P3RDDATA(1)",
          OutTemp       => P3RDDATA_out(1),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(10),
          GlitchData    => P3RDDATA10_GlitchData,
          OutSignalName => "P3RDDATA(10)",
          OutTemp       => P3RDDATA_out(10),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(10),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(11),
          GlitchData    => P3RDDATA11_GlitchData,
          OutSignalName => "P3RDDATA(11)",
          OutTemp       => P3RDDATA_out(11),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(11),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(12),
          GlitchData    => P3RDDATA12_GlitchData,
          OutSignalName => "P3RDDATA(12)",
          OutTemp       => P3RDDATA_out(12),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(12),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(13),
          GlitchData    => P3RDDATA13_GlitchData,
          OutSignalName => "P3RDDATA(13)",
          OutTemp       => P3RDDATA_out(13),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(13),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(14),
          GlitchData    => P3RDDATA14_GlitchData,
          OutSignalName => "P3RDDATA(14)",
          OutTemp       => P3RDDATA_out(14),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(14),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(15),
          GlitchData    => P3RDDATA15_GlitchData,
          OutSignalName => "P3RDDATA(15)",
          OutTemp       => P3RDDATA_out(15),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(15),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(16),
          GlitchData    => P3RDDATA16_GlitchData,
          OutSignalName => "P3RDDATA(16)",
          OutTemp       => P3RDDATA_out(16),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(16),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(17),
          GlitchData    => P3RDDATA17_GlitchData,
          OutSignalName => "P3RDDATA(17)",
          OutTemp       => P3RDDATA_out(17),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(17),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(18),
          GlitchData    => P3RDDATA18_GlitchData,
          OutSignalName => "P3RDDATA(18)",
          OutTemp       => P3RDDATA_out(18),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(18),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(19),
          GlitchData    => P3RDDATA19_GlitchData,
          OutSignalName => "P3RDDATA(19)",
          OutTemp       => P3RDDATA_out(19),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(19),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(2),
          GlitchData    => P3RDDATA2_GlitchData,
          OutSignalName => "P3RDDATA(2)",
          OutTemp       => P3RDDATA_out(2),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(20),
          GlitchData    => P3RDDATA20_GlitchData,
          OutSignalName => "P3RDDATA(20)",
          OutTemp       => P3RDDATA_out(20),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(20),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(21),
          GlitchData    => P3RDDATA21_GlitchData,
          OutSignalName => "P3RDDATA(21)",
          OutTemp       => P3RDDATA_out(21),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(21),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(22),
          GlitchData    => P3RDDATA22_GlitchData,
          OutSignalName => "P3RDDATA(22)",
          OutTemp       => P3RDDATA_out(22),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(22),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(23),
          GlitchData    => P3RDDATA23_GlitchData,
          OutSignalName => "P3RDDATA(23)",
          OutTemp       => P3RDDATA_out(23),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(23),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(24),
          GlitchData    => P3RDDATA24_GlitchData,
          OutSignalName => "P3RDDATA(24)",
          OutTemp       => P3RDDATA_out(24),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(24),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(25),
          GlitchData    => P3RDDATA25_GlitchData,
          OutSignalName => "P3RDDATA(25)",
          OutTemp       => P3RDDATA_out(25),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(25),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(26),
          GlitchData    => P3RDDATA26_GlitchData,
          OutSignalName => "P3RDDATA(26)",
          OutTemp       => P3RDDATA_out(26),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(26),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(27),
          GlitchData    => P3RDDATA27_GlitchData,
          OutSignalName => "P3RDDATA(27)",
          OutTemp       => P3RDDATA_out(27),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(27),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(28),
          GlitchData    => P3RDDATA28_GlitchData,
          OutSignalName => "P3RDDATA(28)",
          OutTemp       => P3RDDATA_out(28),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(28),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(29),
          GlitchData    => P3RDDATA29_GlitchData,
          OutSignalName => "P3RDDATA(29)",
          OutTemp       => P3RDDATA_out(29),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(29),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(3),
          GlitchData    => P3RDDATA3_GlitchData,
          OutSignalName => "P3RDDATA(3)",
          OutTemp       => P3RDDATA_out(3),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(30),
          GlitchData    => P3RDDATA30_GlitchData,
          OutSignalName => "P3RDDATA(30)",
          OutTemp       => P3RDDATA_out(30),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(30),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(31),
          GlitchData    => P3RDDATA31_GlitchData,
          OutSignalName => "P3RDDATA(31)",
          OutTemp       => P3RDDATA_out(31),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(31),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(4),
          GlitchData    => P3RDDATA4_GlitchData,
          OutSignalName => "P3RDDATA(4)",
          OutTemp       => P3RDDATA_out(4),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(5),
          GlitchData    => P3RDDATA5_GlitchData,
          OutSignalName => "P3RDDATA(5)",
          OutTemp       => P3RDDATA_out(5),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(6),
          GlitchData    => P3RDDATA6_GlitchData,
          OutSignalName => "P3RDDATA(6)",
          OutTemp       => P3RDDATA_out(6),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(7),
          GlitchData    => P3RDDATA7_GlitchData,
          OutSignalName => "P3RDDATA(7)",
          OutTemp       => P3RDDATA_out(7),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(8),
          GlitchData    => P3RDDATA8_GlitchData,
          OutSignalName => "P3RDDATA(8)",
          OutTemp       => P3RDDATA_out(8),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(8),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDDATA(9),
          GlitchData    => P3RDDATA9_GlitchData,
          OutSignalName => "P3RDDATA(9)",
          OutTemp       => P3RDDATA_out(9),
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDDATA(9),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3RDOVERFLOW,
          GlitchData    => P3RDOVERFLOW_GlitchData,
          OutSignalName => "P3RDOVERFLOW",
          OutTemp       => P3RDOVERFLOW_out,
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3RDOVERFLOW,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P3WRUNDERRUN,
          GlitchData    => P3WRUNDERRUN_GlitchData,
          OutSignalName => "P3WRUNDERRUN",
          OutTemp       => P3WRUNDERRUN_out,
          Paths       => (0 => (P3CLK_dly'last_event, tpd_P3CLK_P3WRUNDERRUN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4CMDEMPTY,
          GlitchData    => P4CMDEMPTY_GlitchData,
          OutSignalName => "P4CMDEMPTY",
          OutTemp       => P4CMDEMPTY_out,
          Paths       => (0 => (P4CMDCLK_dly'last_event, tpd_P4CMDCLK_P4CMDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4CMDFULL,
          GlitchData    => P4CMDFULL_GlitchData,
          OutSignalName => "P4CMDFULL",
          OutTemp       => P4CMDFULL_out,
          Paths       => (0 => (P4CMDCLK_dly'last_event, tpd_P4CMDCLK_P4CMDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(0),
          GlitchData    => P4COUNT0_GlitchData,
          OutSignalName => "P4COUNT(0)",
          OutTemp       => P4COUNT_out(0),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(1),
          GlitchData    => P4COUNT1_GlitchData,
          OutSignalName => "P4COUNT(1)",
          OutTemp       => P4COUNT_out(1),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(2),
          GlitchData    => P4COUNT2_GlitchData,
          OutSignalName => "P4COUNT(2)",
          OutTemp       => P4COUNT_out(2),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(3),
          GlitchData    => P4COUNT3_GlitchData,
          OutSignalName => "P4COUNT(3)",
          OutTemp       => P4COUNT_out(3),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(4),
          GlitchData    => P4COUNT4_GlitchData,
          OutSignalName => "P4COUNT(4)",
          OutTemp       => P4COUNT_out(4),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(5),
          GlitchData    => P4COUNT5_GlitchData,
          OutSignalName => "P4COUNT(5)",
          OutTemp       => P4COUNT_out(5),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4COUNT(6),
          GlitchData    => P4COUNT6_GlitchData,
          OutSignalName => "P4COUNT(6)",
          OutTemp       => P4COUNT_out(6),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4COUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4EMPTY,
          GlitchData    => P4EMPTY_GlitchData,
          OutSignalName => "P4EMPTY",
          OutTemp       => P4EMPTY_out,
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4EMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4ERROR,
          GlitchData    => P4ERROR_GlitchData,
          OutSignalName => "P4ERROR",
          OutTemp       => P4ERROR_out,
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4ERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4FULL,
          GlitchData    => P4FULL_GlitchData,
          OutSignalName => "P4FULL",
          OutTemp       => P4FULL_out,
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4FULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(0),
          GlitchData    => P4RDDATA0_GlitchData,
          OutSignalName => "P4RDDATA(0)",
          OutTemp       => P4RDDATA_out(0),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(1),
          GlitchData    => P4RDDATA1_GlitchData,
          OutSignalName => "P4RDDATA(1)",
          OutTemp       => P4RDDATA_out(1),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(10),
          GlitchData    => P4RDDATA10_GlitchData,
          OutSignalName => "P4RDDATA(10)",
          OutTemp       => P4RDDATA_out(10),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(10),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(11),
          GlitchData    => P4RDDATA11_GlitchData,
          OutSignalName => "P4RDDATA(11)",
          OutTemp       => P4RDDATA_out(11),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(11),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(12),
          GlitchData    => P4RDDATA12_GlitchData,
          OutSignalName => "P4RDDATA(12)",
          OutTemp       => P4RDDATA_out(12),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(12),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(13),
          GlitchData    => P4RDDATA13_GlitchData,
          OutSignalName => "P4RDDATA(13)",
          OutTemp       => P4RDDATA_out(13),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(13),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(14),
          GlitchData    => P4RDDATA14_GlitchData,
          OutSignalName => "P4RDDATA(14)",
          OutTemp       => P4RDDATA_out(14),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(14),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(15),
          GlitchData    => P4RDDATA15_GlitchData,
          OutSignalName => "P4RDDATA(15)",
          OutTemp       => P4RDDATA_out(15),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(15),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(16),
          GlitchData    => P4RDDATA16_GlitchData,
          OutSignalName => "P4RDDATA(16)",
          OutTemp       => P4RDDATA_out(16),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(16),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(17),
          GlitchData    => P4RDDATA17_GlitchData,
          OutSignalName => "P4RDDATA(17)",
          OutTemp       => P4RDDATA_out(17),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(17),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(18),
          GlitchData    => P4RDDATA18_GlitchData,
          OutSignalName => "P4RDDATA(18)",
          OutTemp       => P4RDDATA_out(18),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(18),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(19),
          GlitchData    => P4RDDATA19_GlitchData,
          OutSignalName => "P4RDDATA(19)",
          OutTemp       => P4RDDATA_out(19),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(19),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(2),
          GlitchData    => P4RDDATA2_GlitchData,
          OutSignalName => "P4RDDATA(2)",
          OutTemp       => P4RDDATA_out(2),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(20),
          GlitchData    => P4RDDATA20_GlitchData,
          OutSignalName => "P4RDDATA(20)",
          OutTemp       => P4RDDATA_out(20),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(20),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(21),
          GlitchData    => P4RDDATA21_GlitchData,
          OutSignalName => "P4RDDATA(21)",
          OutTemp       => P4RDDATA_out(21),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(21),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(22),
          GlitchData    => P4RDDATA22_GlitchData,
          OutSignalName => "P4RDDATA(22)",
          OutTemp       => P4RDDATA_out(22),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(22),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(23),
          GlitchData    => P4RDDATA23_GlitchData,
          OutSignalName => "P4RDDATA(23)",
          OutTemp       => P4RDDATA_out(23),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(23),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(24),
          GlitchData    => P4RDDATA24_GlitchData,
          OutSignalName => "P4RDDATA(24)",
          OutTemp       => P4RDDATA_out(24),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(24),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(25),
          GlitchData    => P4RDDATA25_GlitchData,
          OutSignalName => "P4RDDATA(25)",
          OutTemp       => P4RDDATA_out(25),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(25),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(26),
          GlitchData    => P4RDDATA26_GlitchData,
          OutSignalName => "P4RDDATA(26)",
          OutTemp       => P4RDDATA_out(26),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(26),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(27),
          GlitchData    => P4RDDATA27_GlitchData,
          OutSignalName => "P4RDDATA(27)",
          OutTemp       => P4RDDATA_out(27),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(27),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(28),
          GlitchData    => P4RDDATA28_GlitchData,
          OutSignalName => "P4RDDATA(28)",
          OutTemp       => P4RDDATA_out(28),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(28),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(29),
          GlitchData    => P4RDDATA29_GlitchData,
          OutSignalName => "P4RDDATA(29)",
          OutTemp       => P4RDDATA_out(29),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(29),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(3),
          GlitchData    => P4RDDATA3_GlitchData,
          OutSignalName => "P4RDDATA(3)",
          OutTemp       => P4RDDATA_out(3),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(30),
          GlitchData    => P4RDDATA30_GlitchData,
          OutSignalName => "P4RDDATA(30)",
          OutTemp       => P4RDDATA_out(30),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(30),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(31),
          GlitchData    => P4RDDATA31_GlitchData,
          OutSignalName => "P4RDDATA(31)",
          OutTemp       => P4RDDATA_out(31),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(31),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(4),
          GlitchData    => P4RDDATA4_GlitchData,
          OutSignalName => "P4RDDATA(4)",
          OutTemp       => P4RDDATA_out(4),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(5),
          GlitchData    => P4RDDATA5_GlitchData,
          OutSignalName => "P4RDDATA(5)",
          OutTemp       => P4RDDATA_out(5),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(6),
          GlitchData    => P4RDDATA6_GlitchData,
          OutSignalName => "P4RDDATA(6)",
          OutTemp       => P4RDDATA_out(6),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(7),
          GlitchData    => P4RDDATA7_GlitchData,
          OutSignalName => "P4RDDATA(7)",
          OutTemp       => P4RDDATA_out(7),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(8),
          GlitchData    => P4RDDATA8_GlitchData,
          OutSignalName => "P4RDDATA(8)",
          OutTemp       => P4RDDATA_out(8),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(8),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDDATA(9),
          GlitchData    => P4RDDATA9_GlitchData,
          OutSignalName => "P4RDDATA(9)",
          OutTemp       => P4RDDATA_out(9),
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDDATA(9),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4RDOVERFLOW,
          GlitchData    => P4RDOVERFLOW_GlitchData,
          OutSignalName => "P4RDOVERFLOW",
          OutTemp       => P4RDOVERFLOW_out,
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4RDOVERFLOW,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P4WRUNDERRUN,
          GlitchData    => P4WRUNDERRUN_GlitchData,
          OutSignalName => "P4WRUNDERRUN",
          OutTemp       => P4WRUNDERRUN_out,
          Paths       => (0 => (P4CLK_dly'last_event, tpd_P4CLK_P4WRUNDERRUN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5CMDEMPTY,
          GlitchData    => P5CMDEMPTY_GlitchData,
          OutSignalName => "P5CMDEMPTY",
          OutTemp       => P5CMDEMPTY_out,
          Paths       => (0 => (P5CMDCLK_dly'last_event, tpd_P5CMDCLK_P5CMDEMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5CMDFULL,
          GlitchData    => P5CMDFULL_GlitchData,
          OutSignalName => "P5CMDFULL",
          OutTemp       => P5CMDFULL_out,
          Paths       => (0 => (P5CMDCLK_dly'last_event, tpd_P5CMDCLK_P5CMDFULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(0),
          GlitchData    => P5COUNT0_GlitchData,
          OutSignalName => "P5COUNT(0)",
          OutTemp       => P5COUNT_out(0),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(1),
          GlitchData    => P5COUNT1_GlitchData,
          OutSignalName => "P5COUNT(1)",
          OutTemp       => P5COUNT_out(1),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(2),
          GlitchData    => P5COUNT2_GlitchData,
          OutSignalName => "P5COUNT(2)",
          OutTemp       => P5COUNT_out(2),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(3),
          GlitchData    => P5COUNT3_GlitchData,
          OutSignalName => "P5COUNT(3)",
          OutTemp       => P5COUNT_out(3),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(4),
          GlitchData    => P5COUNT4_GlitchData,
          OutSignalName => "P5COUNT(4)",
          OutTemp       => P5COUNT_out(4),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(5),
          GlitchData    => P5COUNT5_GlitchData,
          OutSignalName => "P5COUNT(5)",
          OutTemp       => P5COUNT_out(5),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5COUNT(6),
          GlitchData    => P5COUNT6_GlitchData,
          OutSignalName => "P5COUNT(6)",
          OutTemp       => P5COUNT_out(6),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5COUNT(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5EMPTY,
          GlitchData    => P5EMPTY_GlitchData,
          OutSignalName => "P5EMPTY",
          OutTemp       => P5EMPTY_out,
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5EMPTY,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5ERROR,
          GlitchData    => P5ERROR_GlitchData,
          OutSignalName => "P5ERROR",
          OutTemp       => P5ERROR_out,
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5ERROR,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5FULL,
          GlitchData    => P5FULL_GlitchData,
          OutSignalName => "P5FULL",
          OutTemp       => P5FULL_out,
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5FULL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(0),
          GlitchData    => P5RDDATA0_GlitchData,
          OutSignalName => "P5RDDATA(0)",
          OutTemp       => P5RDDATA_out(0),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(1),
          GlitchData    => P5RDDATA1_GlitchData,
          OutSignalName => "P5RDDATA(1)",
          OutTemp       => P5RDDATA_out(1),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(10),
          GlitchData    => P5RDDATA10_GlitchData,
          OutSignalName => "P5RDDATA(10)",
          OutTemp       => P5RDDATA_out(10),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(10),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(11),
          GlitchData    => P5RDDATA11_GlitchData,
          OutSignalName => "P5RDDATA(11)",
          OutTemp       => P5RDDATA_out(11),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(11),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(12),
          GlitchData    => P5RDDATA12_GlitchData,
          OutSignalName => "P5RDDATA(12)",
          OutTemp       => P5RDDATA_out(12),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(12),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(13),
          GlitchData    => P5RDDATA13_GlitchData,
          OutSignalName => "P5RDDATA(13)",
          OutTemp       => P5RDDATA_out(13),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(13),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(14),
          GlitchData    => P5RDDATA14_GlitchData,
          OutSignalName => "P5RDDATA(14)",
          OutTemp       => P5RDDATA_out(14),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(14),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(15),
          GlitchData    => P5RDDATA15_GlitchData,
          OutSignalName => "P5RDDATA(15)",
          OutTemp       => P5RDDATA_out(15),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(15),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(16),
          GlitchData    => P5RDDATA16_GlitchData,
          OutSignalName => "P5RDDATA(16)",
          OutTemp       => P5RDDATA_out(16),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(16),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(17),
          GlitchData    => P5RDDATA17_GlitchData,
          OutSignalName => "P5RDDATA(17)",
          OutTemp       => P5RDDATA_out(17),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(17),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(18),
          GlitchData    => P5RDDATA18_GlitchData,
          OutSignalName => "P5RDDATA(18)",
          OutTemp       => P5RDDATA_out(18),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(18),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(19),
          GlitchData    => P5RDDATA19_GlitchData,
          OutSignalName => "P5RDDATA(19)",
          OutTemp       => P5RDDATA_out(19),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(19),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(2),
          GlitchData    => P5RDDATA2_GlitchData,
          OutSignalName => "P5RDDATA(2)",
          OutTemp       => P5RDDATA_out(2),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(20),
          GlitchData    => P5RDDATA20_GlitchData,
          OutSignalName => "P5RDDATA(20)",
          OutTemp       => P5RDDATA_out(20),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(20),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(21),
          GlitchData    => P5RDDATA21_GlitchData,
          OutSignalName => "P5RDDATA(21)",
          OutTemp       => P5RDDATA_out(21),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(21),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(22),
          GlitchData    => P5RDDATA22_GlitchData,
          OutSignalName => "P5RDDATA(22)",
          OutTemp       => P5RDDATA_out(22),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(22),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(23),
          GlitchData    => P5RDDATA23_GlitchData,
          OutSignalName => "P5RDDATA(23)",
          OutTemp       => P5RDDATA_out(23),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(23),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(24),
          GlitchData    => P5RDDATA24_GlitchData,
          OutSignalName => "P5RDDATA(24)",
          OutTemp       => P5RDDATA_out(24),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(24),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(25),
          GlitchData    => P5RDDATA25_GlitchData,
          OutSignalName => "P5RDDATA(25)",
          OutTemp       => P5RDDATA_out(25),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(25),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(26),
          GlitchData    => P5RDDATA26_GlitchData,
          OutSignalName => "P5RDDATA(26)",
          OutTemp       => P5RDDATA_out(26),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(26),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(27),
          GlitchData    => P5RDDATA27_GlitchData,
          OutSignalName => "P5RDDATA(27)",
          OutTemp       => P5RDDATA_out(27),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(27),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(28),
          GlitchData    => P5RDDATA28_GlitchData,
          OutSignalName => "P5RDDATA(28)",
          OutTemp       => P5RDDATA_out(28),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(28),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(29),
          GlitchData    => P5RDDATA29_GlitchData,
          OutSignalName => "P5RDDATA(29)",
          OutTemp       => P5RDDATA_out(29),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(29),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(3),
          GlitchData    => P5RDDATA3_GlitchData,
          OutSignalName => "P5RDDATA(3)",
          OutTemp       => P5RDDATA_out(3),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(30),
          GlitchData    => P5RDDATA30_GlitchData,
          OutSignalName => "P5RDDATA(30)",
          OutTemp       => P5RDDATA_out(30),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(30),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(31),
          GlitchData    => P5RDDATA31_GlitchData,
          OutSignalName => "P5RDDATA(31)",
          OutTemp       => P5RDDATA_out(31),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(31),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(4),
          GlitchData    => P5RDDATA4_GlitchData,
          OutSignalName => "P5RDDATA(4)",
          OutTemp       => P5RDDATA_out(4),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(5),
          GlitchData    => P5RDDATA5_GlitchData,
          OutSignalName => "P5RDDATA(5)",
          OutTemp       => P5RDDATA_out(5),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(6),
          GlitchData    => P5RDDATA6_GlitchData,
          OutSignalName => "P5RDDATA(6)",
          OutTemp       => P5RDDATA_out(6),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(7),
          GlitchData    => P5RDDATA7_GlitchData,
          OutSignalName => "P5RDDATA(7)",
          OutTemp       => P5RDDATA_out(7),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(8),
          GlitchData    => P5RDDATA8_GlitchData,
          OutSignalName => "P5RDDATA(8)",
          OutTemp       => P5RDDATA_out(8),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(8),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDDATA(9),
          GlitchData    => P5RDDATA9_GlitchData,
          OutSignalName => "P5RDDATA(9)",
          OutTemp       => P5RDDATA_out(9),
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDDATA(9),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5RDOVERFLOW,
          GlitchData    => P5RDOVERFLOW_GlitchData,
          OutSignalName => "P5RDOVERFLOW",
          OutTemp       => P5RDOVERFLOW_out,
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5RDOVERFLOW,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => P5WRUNDERRUN,
          GlitchData    => P5WRUNDERRUN_GlitchData,
          OutSignalName => "P5WRUNDERRUN",
          OutTemp       => P5WRUNDERRUN_out,
          Paths       => (0 => (P5CLK_dly'last_event, tpd_P5CLK_P5WRUNDERRUN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => SELFREFRESHMODE,
          GlitchData    => SELFREFRESHMODE_GlitchData,
          OutSignalName => "SELFREFRESHMODE",
          OutTemp       => SELFREFRESHMODE_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_SELFREFRESHMODE(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => SELFREFRESHMODE,
          GlitchData    => SELFREFRESHMODE_GlitchData,
          OutSignalName => "SELFREFRESHMODE",
          OutTemp       => SELFREFRESHMODE_out,
          Paths       => (0 => (PLLCLK_dly'last_event, tpd_PLLCLK_SELFREFRESHMODE(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UOCALSTART,
          GlitchData    => UOCALSTART_GlitchData,
          OutSignalName => "UOCALSTART",
          OutTemp       => UOCALSTART_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UOCALSTART,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UOCMDREADYIN,
          GlitchData    => UOCMDREADYIN_GlitchData,
          OutSignalName => "UOCMDREADYIN",
          OutTemp       => UOCMDREADYIN_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UOCMDREADYIN,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(0),
          GlitchData    => UODATA0_GlitchData,
          OutSignalName => "UODATA(0)",
          OutTemp       => UODATA_out(0),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(0),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(1),
          GlitchData    => UODATA1_GlitchData,
          OutSignalName => "UODATA(1)",
          OutTemp       => UODATA_out(1),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(1),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(2),
          GlitchData    => UODATA2_GlitchData,
          OutSignalName => "UODATA(2)",
          OutTemp       => UODATA_out(2),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(2),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(3),
          GlitchData    => UODATA3_GlitchData,
          OutSignalName => "UODATA(3)",
          OutTemp       => UODATA_out(3),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(3),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(4),
          GlitchData    => UODATA4_GlitchData,
          OutSignalName => "UODATA(4)",
          OutTemp       => UODATA_out(4),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(4),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(5),
          GlitchData    => UODATA5_GlitchData,
          OutSignalName => "UODATA(5)",
          OutTemp       => UODATA_out(5),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(5),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(6),
          GlitchData    => UODATA6_GlitchData,
          OutSignalName => "UODATA(6)",
          OutTemp       => UODATA_out(6),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(6),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATA(7),
          GlitchData    => UODATA7_GlitchData,
          OutSignalName => "UODATA(7)",
          OutTemp       => UODATA_out(7),
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATA(7),TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODATAVALID,
          GlitchData    => UODATAVALID_GlitchData,
          OutSignalName => "UODATAVALID",
          OutTemp       => UODATAVALID_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODATAVALID,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UODONECAL,
          GlitchData    => UODONECAL_GlitchData,
          OutSignalName => "UODONECAL",
          OutTemp       => UODONECAL_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UODONECAL,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UOREFRSHFLAG,
          GlitchData    => UOREFRSHFLAG_GlitchData,
          OutSignalName => "UOREFRSHFLAG",
          OutTemp       => UOREFRSHFLAG_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UOREFRSHFLAG,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPathDelay01
        (
          OutSignal     => UOSDO,
          GlitchData    => UOSDO_GlitchData,
          OutSignalName => "UOSDO",
          OutTemp       => UOSDO_out,
          Paths       => (0 => (UICLK_dly'last_event, tpd_UICLK_UOSDO,TRUE)),
          Mode          => VitalTransport,
          Xon           => false,
          MsgOn          => false,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P0CMDCLK,
          PeriodData     => PInfo_P0CMDCLK,
          TestSignal     => P0CMDCLK_dly,
          TestSignalName => "P0CMDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P0CMDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P0RDCLK,
          PeriodData     => PInfo_P0RDCLK,
          TestSignal     => P0RDCLK_dly,
          TestSignalName => "P0RDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P0RDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P0WRCLK,
          PeriodData     => PInfo_P0WRCLK,
          TestSignal     => P0WRCLK_dly,
          TestSignalName => "P0WRCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P0WRCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P1CMDCLK,
          PeriodData     => PInfo_P1CMDCLK,
          TestSignal     => P1CMDCLK_dly,
          TestSignalName => "P1CMDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P1CMDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P1RDCLK,
          PeriodData     => PInfo_P1RDCLK,
          TestSignal     => P1RDCLK_dly,
          TestSignalName => "P1RDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P1RDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P1WRCLK,
          PeriodData     => PInfo_P1WRCLK,
          TestSignal     => P1WRCLK_dly,
          TestSignalName => "P1WRCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P1WRCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P2CLK,
          PeriodData     => PInfo_P2CLK,
          TestSignal     => P2CLK_dly,
          TestSignalName => "P2CLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P2CLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P2CMDCLK,
          PeriodData     => PInfo_P2CMDCLK,
          TestSignal     => P2CMDCLK_dly,
          TestSignalName => "P2CMDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P2CMDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P3CLK,
          PeriodData     => PInfo_P3CLK,
          TestSignal     => P3CLK_dly,
          TestSignalName => "P3CLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P3CLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P3CMDCLK,
          PeriodData     => PInfo_P3CMDCLK,
          TestSignal     => P3CMDCLK_dly,
          TestSignalName => "P3CMDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P3CMDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P4CLK,
          PeriodData     => PInfo_P4CLK,
          TestSignal     => P4CLK_dly,
          TestSignalName => "P4CLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P4CLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P4CMDCLK,
          PeriodData     => PInfo_P4CMDCLK,
          TestSignal     => P4CMDCLK_dly,
          TestSignalName => "P4CMDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P4CMDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P5CLK,
          PeriodData     => PInfo_P5CLK,
          TestSignal     => P5CLK_dly,
          TestSignalName => "P5CLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P5CLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_P5CMDCLK,
          PeriodData     => PInfo_P5CMDCLK,
          TestSignal     => P5CMDCLK_dly,
          TestSignalName => "P5CMDCLK",
          TestDelay      => 0 ps,
          Period         => tperiod_P5CMDCLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_PLLCLK(0),
          PeriodData     => PInfo_PLLCLK,
          TestSignal     => PLLCLK_dly(0),
          TestSignalName => "PLLCLK(0)",
          TestDelay      => 0 ps,
          Period         => tperiod_PLLCLK_posedge(0),
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
         VitalPeriodPulseCheck
        (
          Violation      => Pviol_PLLCLK(1),
          PeriodData     => PInfo_PLLCLK,
          TestSignal     => PLLCLK_dly(1),
          TestSignalName => "PLLCLK(1)",
          TestDelay      => 0 ps,
          Period         => tperiod_PLLCLK_posedge(1),
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );

        VitalPeriodPulseCheck
        (
          Violation      => Pviol_SYSRST,
          PeriodData     => PInfo_SYSRST,
          TestSignal     => SYSRST_dly,
          TestSignalName => "SYSRST",
          TestDelay      => 0 ps,
          Period         => tperiod_SYSRST_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
        VitalPeriodPulseCheck
        (
          Violation      => Pviol_UICLK,
          PeriodData     => PInfo_UICLK,
          TestSignal     => UICLK_dly,
          TestSignalName => "UICLK",
          TestDelay      => 0 ps,
          Period         => tperiod_UICLK_posedge,
          PulseWidthHigh => 0 ps,
          PulseWidthLow  => 0 ps,
          CheckEnabled   => TRUE,
          HeaderMsg      => InstancePath & "/X_MCB",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity    => WARNING
        );
      wait on
        ADDR_out,
        BA_out,
        CAS_out,
        CKE_out,
        DQIOWEN0_out,
        DQON_out,
        DQOP_out,
        DQSIOWEN90N_out,
        DQSIOWEN90P_out,
        IOIDRPADDR_out,
        IOIDRPADD_out,
        IOIDRPBROADCAST_out,
        IOIDRPCLK_out,
        IOIDRPCS_out,
        IOIDRPSDO_out,
        IOIDRPTRAIN_out,
        IOIDRPUPDATE_out,
        LDMN_out,
        LDMP_out,
        ODT_out,
        P0CMDEMPTY_out,
        P0CMDFULL_out,
        P0RDCOUNT_out,
        P0RDDATA_out,
        P0RDEMPTY_out,
        P0RDERROR_out,
        P0RDFULL_out,
        P0RDOVERFLOW_out,
        P0WRCOUNT_out,
        P0WREMPTY_out,
        P0WRERROR_out,
        P0WRFULL_out,
        P0WRUNDERRUN_out,
        P1CMDEMPTY_out,
        P1CMDFULL_out,
        P1RDCOUNT_out,
        P1RDDATA_out,
        P1RDEMPTY_out,
        P1RDERROR_out,
        P1RDFULL_out,
        P1RDOVERFLOW_out,
        P1WRCOUNT_out,
        P1WREMPTY_out,
        P1WRERROR_out,
        P1WRFULL_out,
        P1WRUNDERRUN_out,
        P2CMDEMPTY_out,
        P2CMDFULL_out,
        P2COUNT_out,
        P2EMPTY_out,
        P2ERROR_out,
        P2FULL_out,
        P2RDDATA_out,
        P2RDOVERFLOW_out,
        P2WRUNDERRUN_out,
        P3CMDEMPTY_out,
        P3CMDFULL_out,
        P3COUNT_out,
        P3EMPTY_out,
        P3ERROR_out,
        P3FULL_out,
        P3RDDATA_out,
        P3RDOVERFLOW_out,
        P3WRUNDERRUN_out,
        P4CMDEMPTY_out,
        P4CMDFULL_out,
        P4COUNT_out,
        P4EMPTY_out,
        P4ERROR_out,
        P4FULL_out,
        P4RDDATA_out,
        P4RDOVERFLOW_out,
        P4WRUNDERRUN_out,
        P5CMDEMPTY_out,
        P5CMDFULL_out,
        P5COUNT_out,
        P5EMPTY_out,
        P5ERROR_out,
        P5FULL_out,
        P5RDDATA_out,
        P5RDOVERFLOW_out,
        P5WRUNDERRUN_out,
        RAS_out,
        RST_out,
        SELFREFRESHMODE_out,
        STATUS_out,
        UDMN_out,
        UDMP_out,
        UOCALSTART_out,
        UOCMDREADYIN_out,
        UODATAVALID_out,
        UODATA_out,
        UODONECAL_out,
        UOREFRSHFLAG_out,
        UOSDO_out,
        WE_out,
        IOIDRPSDI_UICLK_dly,
        P0ARBEN_PLLCLK_dly,
        P0CMDBA_P0CMDCLK_dly,
        P0CMDBL_P0CMDCLK_dly,
        P0CMDCA_P0CMDCLK_dly,
        P0CMDEN_P0CMDCLK_dly,
        P0CMDINSTR_P0CMDCLK_dly,
        P0CMDRA_P0CMDCLK_dly,
        P0RDEN_P0RDCLK_dly,
        P0RWRMASK_P0WRCLK_dly,
        P0WRDATA_P0WRCLK_dly,
        P0WREN_P0WRCLK_dly,
        P1ARBEN_PLLCLK_dly,
        P1CMDBA_P1CMDCLK_dly,
        P1CMDBL_P1CMDCLK_dly,
        P1CMDCA_P1CMDCLK_dly,
        P1CMDEN_P1CMDCLK_dly,
        P1CMDINSTR_P1CMDCLK_dly,
        P1CMDRA_P1CMDCLK_dly,
        P1RDEN_P1RDCLK_dly,
        P1RWRMASK_P1WRCLK_dly,
        P1WRDATA_P1WRCLK_dly,
        P1WREN_P1WRCLK_dly,
        P2ARBEN_PLLCLK_dly,
        P2CMDBA_P2CMDCLK_dly,
        P2CMDBL_P2CMDCLK_dly,
        P2CMDCA_P2CMDCLK_dly,
        P2CMDEN_P2CMDCLK_dly,
        P2CMDINSTR_P2CMDCLK_dly,
        P2CMDRA_P2CMDCLK_dly,
        P2EN_P2CLK_dly,
        P2WRDATA_P2CLK_dly,
        P2WRMASK_P2CLK_dly,
        P3ARBEN_PLLCLK_dly,
        P3CMDBA_P3CMDCLK_dly,
        P3CMDBL_P3CMDCLK_dly,
        P3CMDCA_P3CMDCLK_dly,
        P3CMDEN_P3CMDCLK_dly,
        P3CMDINSTR_P3CMDCLK_dly,
        P3CMDRA_P3CMDCLK_dly,
        P3EN_P3CLK_dly,
        P3WRDATA_P3CLK_dly,
        P3WRMASK_P3CLK_dly,
        P4ARBEN_PLLCLK_dly,
        P4CMDBA_P4CMDCLK_dly,
        P4CMDBL_P4CMDCLK_dly,
        P4CMDCA_P4CMDCLK_dly,
        P4CMDEN_P4CMDCLK_dly,
        P4CMDINSTR_P4CMDCLK_dly,
        P4CMDRA_P4CMDCLK_dly,
        P4EN_P4CLK_dly,
        P4WRDATA_P4CLK_dly,
        P4WRMASK_P4CLK_dly,
        P5ARBEN_PLLCLK_dly,
        P5CMDBA_P5CMDCLK_dly,
        P5CMDBL_P5CMDCLK_dly,
        P5CMDCA_P5CMDCLK_dly,
        P5CMDEN_P5CMDCLK_dly,
        P5CMDINSTR_P5CMDCLK_dly,
        P5CMDRA_P5CMDCLK_dly,
        P5EN_P5CLK_dly,
        P5WRDATA_P5CLK_dly,
        P5WRMASK_P5CLK_dly,
        PLLCE_PLLCLK_dly,
        PLLLOCK_PLLCLK_dly,
        RECAL_PLLCLK_dly,
        SELFREFRESHENTER_PLLCLK_dly,
        UIADDR_UICLK_dly,
        UIADD_UICLK_dly,
        UIBROADCAST_UICLK_dly,
        UICMDEN_UICLK_dly,
        UICMDIN_UICLK_dly,
        UICMD_UICLK_dly,
        UICS_UICLK_dly,
        UIDONECAL_UICLK_dly,
        UIDQCOUNT_UICLK_dly,
        UIDQLOWERDEC_UICLK_dly,
        UIDQLOWERINC_UICLK_dly,
        UIDQUPPERDEC_UICLK_dly,
        UIDQUPPERINC_UICLK_dly,
        UIDRPUPDATE_UICLK_dly,
        UILDQSDEC_UICLK_dly,
        UILDQSINC_UICLK_dly,
        UIREAD_UICLK_dly,
        UISDI_UICLK_dly,
        UIUDQSDEC_UICLK_dly,
        UIUDQSINC_UICLK_dly;
    end process TIMING;
    ADDR <= ADDR_out;
    BA <= BA_out;
    CAS <= CAS_out;
    CKE <= CKE_out;
    DQON <= DQON_out;
    DQOP <= DQOP_out;
    IOIDRPTRAIN <= IOIDRPTRAIN_out;
    LDMN <= LDMN_out;
    LDMP <= LDMP_out;
    ODT <= ODT_out;
    RAS <= RAS_out;
    RST <= RST_out;
    STATUS <= STATUS_out;
    UDMN <= UDMN_out;
    UDMP <= UDMP_out;
    WE <= WE_out;
  end X_MCB_V;
