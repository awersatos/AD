*=======================================================
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.
*/////////////////////////////////////////////////////////////////////
* Legal Notice:
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice.
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND"
*////////////////////////////////////////////////////////////////////
* For more information, and our latest models,
* please visit the models section of our website at
*       http://www.national.com/models/
*////////////////////////////////////////////////////////////////////
*
* Rev 1.8 (2008/11/03) PG - Connected Q13/14 Substrate directly to VEE, removed R100.
* Rev 1.7 (2008/07/28) PG - Release Rev.
*
*
*
* PARAMETERS NOT MODELLED:
* -Distortion
* -Noise
* -CMVR (Common Mode Voltage Range)
* -Common-mode control loop behavior (Vcm_ref to output)
* -Temperature effects
* -Differential Offset Voltage
* -Gain/ Phase Balance Error
* -Common Mode Gain (input to output)
* -PSRR (Common Mode and Differential Mode)
* Vcm_REF input current when clamped (> 1.9V, < 0.7V)
*********
* PARAMETERS MODELED LOOSELY:
* -Output voltage range
* -Vcm_REF voltage range
* -Undriven input response (single ended input drive)
* -Input common mode with source resistance
* -output response with Vout > 800mVpp
*
* PINOUT ORDER +IN -IN V+ V- +OUT -OUT VCM
* PINOUT ORDER  16  5  12 1    8   13   10

.subckt LMH6555 VINP VINN VCC VEE VOUTP VOUTN VCMREFIN

D2 a130 a0177 DIODEnoisy
D3 a111 a117 DIODEnoisy
G1 a071 VEE a081 VCMREF 10m
G0 a138 VEE a081 VCMREF 10m
E8 a0141 VEE a075 VEE 1.0
E0 a073 0 a0101 0 1.0
E2 a138 a071 a0162 0 1000
C9 a081 VEE 10p
C5 a0162 0 101f
C1 a0101 0 26.5p
Q13 VCC a138 op VEE NPNXTR
Q14 VCC a071 on VEE NPNXTR
V15 VCC a76 0
V5 a0152 0 0
V4 a0113 0 0
V1 a130 a111 0
V16 a177 VEE 0
I12 a0177 a117 0m
I5 VCC VCMREF 12u
I46 a76 a177 46.7m
F11 VCC a130 V15 .1801
F12 VCC a111 V15 .1801
F16 op VEE V16 .55675
F17 on VEE V16 .55675
F4 VCC a111 V4 1.0
F5 VCC a130 V5 1.0
F0 0 a0101 V1 .1866
R44 VINP a0177 40.32
R43 a117 VINN 40.32
R42 on a0177 440
R41 a117 op 440
R56 a081 a0141 1K
R50 on VOUTN 50
RTM a0101 0 1K
RGM a117 VEE 32
R26 a0152 0 320
R25 a0113 0 320
R15 op a075 100
R16 a075 on 100
RGP a0177 VEE 32
R49 op VOUTP 50
R51 a073 a0162 1K
DCOPN a2001 op DIODEideal
VCOPN VEE a2001 -1
DCONN a2003 on DIODEideal
VCONN VEE a2003 -1
VCVCMP VCC a2004 2.2
DCVCMP VCMREF a2004 DIODEideal
DCVCMN a2005 VCMREF DIODEideal
VCVCMN VEE a2005 -1.3
RVCM VCMREF VCMREFIN 0.1

* Models
.model DIODEideal d(tnom=25.0 is=1e-18)
.model DIODEnoisy d(tnom=25.0 is=1e-18 af=2.0 kf=80e-12)
.model NPNXTR npn(tnom=25.0 is=14.42e-18 bf=300
+  vaf=200.0 rb=57.00 re=3.000
+  rc=7.000  cje=206.3e-15  cjc=81.45e-15
+  kf=480.0e-12 af=2.000)


.ends LMH6555

