* BEGIN MODEL LMH6321
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.
*/////////////////////////////////////////////////////////////////////
* Legal Notice:
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice.
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND"
*////////////////////////////////////////////////////////////////////
* Rev 1.01
* Fixed IKF typo in NPN model in line 116 - 5/23/08 PG
*
*

* PINOUT ORDER IN V+ V- OUT
* PINOUT ORDER 3  77 44  6

* BEGIN NOTES
* MODEL DOES NOT HAVE PROGRAMMABLE CURRENT LIMIT
* MODEL FEATURES ARE
* GAIN
* SLEW
* SWING
* VOLTAGE NOISE
* CURRENT NOISE
* INPUT BIAS CURRENT
* POWER SUPPLY REJECTION
* QUIESCENT CURRENT
* END NOTES

.SUBCKT LMH6321 3 77 44 6
R4 80 85 50
Q4 44 85 87 7 QP 4
Q5 88 88 86 7 QP 4
R5 92 77 400
Q9 90 92 92 7 QP 4
R6 93 77 270
Q10 90 94 93 7 QP 2
R7 95 77 400
C1 95 90 0.5E-12
Q11 89 96 96 4 Q 8
R12 102 84 30
Q14 44 103 94 7 QP
Q15 44 104 105 7 QP 12
R13 105 85 50
R15 90 100 50
R16 89 104 150
R17 91 108 15
R1 82 79 1
R18 88 110 15
R19 111 109 65
Q21 44 114 99 7 QP
Q22 114 114 115 7 QP
R22 44 114 1600
Q23 77 99 116 4 Q
R23 44 116 1600
Q24 103 117 99 4 Q
Q25 117 117 115 4 Q
I1 77 117 160E-6
Q26 118 118 113 4 Q
Q27 77 118 94 4 Q
R24 118 77 1200
R25 93 119 100
Q6 89 89 88 7 QP 4
R26 98 120 100
Q28 90 121 6 4 QNI 8
R29 82 121 50
Q29 89 122 6 7 QPI 8
R31 83 122 50
Q3 77 84 86 4 Q 4
R32 6 82 1.1
R33 81 83 1
Q1 77 78 79 4 QNO 7.5
R2 83 6 1.1
R3 78 84 150
M2 123 106 119 119 M3N
R35 123 119 3
R14 85 106 30
Q16 77 107 106 4 Q 12
Q17 77 107 108 4 Q 4
Q18 44 109 102 7 QP 12
Q19 44 109 110 7 QP 4
Q30 124 125 119 4 Q
R36 123 125 100
D2 106 124 DD
R38 126 120 3
R8 44 96 400
R9 44 97 400
C2 89 97 0.5E-12
R10 44 98 202
Q12 89 99 98 4 Q 2
Q13 77 100 101 4 Q 12
R11 84 101 50
M3 126 102 120 120 M3P
Q2 44 80 81 7 QPO 8.6
Q31 127 128 120 7 QP
R39 126 128 100
D3 127 102 DD
R20 107 111 65
R21 111 112 65
Q20 103 103 113 7 QP
Q7 90 90 91 4 Q 4
Q8 91 91 87 4 Q 4
V4 3 112 -16E-3
E1 7 0 77 0 1
E2 4 0 44 0 1
R40 0 7 1E12
R41 0 4 1E12
R42 0 4 1E12
R43 0 7 1E12
.MODEL QNI NPN
.MODEL QPI PNP
.MODEL Q NPN  IS=1.76E-16 BF=170 NF=1 VAF=335 IKF=0.08 ISE=6E-16 NE=1.6
+ BR=0.36 NR=1 VAR=3 IKR=6.88E-05 ISC=2.4E-15 NC=1 RB=113.1 IRB=1.23E-4
+ RBM=18.4 RE=1.19 RC=19.6 XTI=2 EG=1.17 XTB=1.2 AF=1 KF=1E-18
+ TF=4.20E-11 XTF=118 ITF=1.6E-2 VTF=0.42 PTF=45 TR=5E-09 CJE=4.8E-13
+ VJE=0.94 MJE=0.42 FC=0.5 CJC=2.75E-13 VJC=0.75 MJC=0.42 CJS=1.01E-12
+ VJS=0.67 MJS=0.322
.MODEL QP PNP IS=2.00E-16 BF=80 NF=1 VAF=118 IKF=0.02 ISE=8E-16 NE=1.65
+ BR=0.14 NR=1 VAR=2 IKR=1E-4 ISC=5.60E-15 NC=1 RB=44.8 IRB=1.5E-4
+ RBM=13.8 RE=1.88 RC=35 XTI=2 EG=1.17 XTB=1.2 AF=1 KF=1E-18 TF=9.40E-11
+ XTF=36.8 ITF=1.34E-2 VTF=1.14 PTF=45 TR=5E-09 CJE=4.32E-13 VJE=0.95
+ MJE=0.38 FC=0.5 CJC=4.84E-13 VJC=0.7 MJC=0.47 CJS=1.42E-12 VJS=0.8
+ MJS=0.23
.MODEL QNO NPN IS=1.41E-15 BF=170 NF=1 VAF=335 IKF=0.64 ISE=4.8E-15 NE=1.6
+ BR=0.36 NR=1 VAR=3 IKR=5.5E-4 ISC=1.92E-14 NC=1 RB=18.3 IRB=9.41E-4
+ RBM=4.14 RE=0.586 RC=8.98 XTI=2 EG=1.17 XTB=1.2 AF=1 KF=1E-18
+ TF=4.2E-11 XTF=118 ITF=1.28E-1 VTF=0.42 PTF=45 TR=5E-09 CJE=3.84E-12
+ VJE=0.94 MJE=0.42 FC=0.5 CJC=1.54E-12 VJC=0.75 MJC=0.42 CJS=3.07E-12
+ VJS=0.67 MJS=0.322
.MODEL QPO PNP IS=1.60E-15 BF=80 NF=1 VAF=118 IKF=0.16 ISE=6.40E-15 NE=1.65
+ BR=0.14 NR=1 VAR=2 IKR=8E-4 ISC=4.48E-14 NC=1 RB=8.48 IRB=1.14E-3
+ RBM=3.55 RE=0.672 RC=18.4 XTI=2 EG=1.17 XTB=1.2 AF=1 KF=1E-18 TF=9.40E-11
+ XTF=36.8 ITF=1.075E-1 VTF=1.14 PTF=45 TR=5E-09 CJE=3.46E-12 VJE=0.95
+ MJE=0.38 FC=0.5 CJC=2.72E-12 VJC=0.7 MJC=0.47 CJS=3.75E-12 VJS=0.8
+ MJS=0.23
.MODEL M3N NMOS VTO=2 KP=0.085 RD=0.1 RS=0.05 IS=1E-18  CGSO=8E-8
+ CGDO=2E-8
.MODEL M3P PMOS VTO=-2 KP=0.085 RD=0.1 RS=0.05 IS=1E-18  CGSO=8E-8
+ CGDO=2E-8
.MODEL DD D RS=1E3 CJO=12E-15 IS=1.72E-17
.ENDS
* END MODEL LMH6321

