*MAC15A8 MCE 2-27-96
*600V 15A pkg:TO-220 2,3,1
.SUBCKT MAC15A8   1  2  3
*     TERMINALS: MT2 G MT1
QN1  5 4 3  NOUT OFF
QN2 11 6 7  NOUT OFF
QP1 6 11 3  POUT OFF
QP2  4 5 7  POUT OFF
DF  4  5  DZ OFF
DR  6 11  DZ OFF
RF  4 6  60MEG
RT2 1 7  18.8M
RH  7 6  87.5
RGP 8 3  23.1
RG  2 8  11.5
RS  8 4  102
DN  9 2  DIN OFF
RN  9 3  41.6
GNN  6 7 9 3 15.2M
GNP  4 5 9 3 18.1M
DP 2 10  DIP OFF
RP 10 3  29.5
GP  7 6 10 3 10.3M
.MODEL DIN  D (IS=45.8F)
.MODEL DIP  D (IS=45.8F N=1.2)
.MODEL DZ   D (IS=45.8F N=1.5 IBV=10U BV=600)
.MODEL POUT PNP (IS=45.8F BF=5 CJE=4.02N TF=38.2U)
.MODEL NOUT NPN (IS=45.8F BF=20 CJE=4.02N CJC=804P TF=2.55U)
.ENDS MAC15A8