`resetall
`timescale 1 ns / 1 ps
`celldefine
module PVTIOCTRL (UPDATE);
  input UPDATE;

endmodule
`endcelldefine
