--------------------------------------------------------------------
--       Actel IGLOO Vital Library
--       NAME: igloo.vhd
--       DATE: September 4, 2007
---------------------------------------------------------------------/

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;

package COMPONENTS is

constant DefaultTimingChecksOn : Boolean := True;
constant DefaultXGenerationOn  : Boolean := False;
constant DefaultXon            : Boolean := False;
constant DefaultMsgOn          : Boolean := True;

component DYNCCC
   generic(
      VCOFREQUENCY      :  Real    := 0.0;
      f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

      TimingChecksOn    :  Boolean := True;
      InstancePath      :  STRING  := "*";
      Xon               :  Boolean := False;
      MsgOn             :  Boolean := True;

      tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKC         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SDIN         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SCLK         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SSHIFT       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SUPDATE      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_MODE         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

      tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );

      tpd_SCLK_SDOUT    : VitalDelayType01  := ( 0.100 ns, 0.100 ns );

      tsetup_SSHIFT_SCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_SSHIFT_SCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_negedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_SDIN_SCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_SDIN_SCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_negedge_posedge    : VitalDelayType := 0.000 ns;

      tpw_SUPDATE_posedge                : VitalDelayType := 0.000 ns;
      tpw_SUPDATE_negedge                : VitalDelayType := 0.000 ns;
      tpw_SCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_SCLK_negedge                   : VitalDelayType := 0.000 ns

      ); 

   port (
          CLKA         : in    std_ulogic;
          EXTFB        : in    std_ulogic;
          POWERDOWN    : in    std_ulogic;
          CLKB         : in    std_ulogic;
          CLKC         : in    std_ulogic;
          SDIN         : in    std_ulogic;
          SCLK         : in    std_ulogic;
          SSHIFT       : in    std_ulogic;
          SUPDATE      : in    std_ulogic;
          MODE         : in    std_ulogic;
          OADIV0       : in    std_ulogic;
          OADIV1       : in    std_ulogic;
          OADIV2       : in    std_ulogic;
          OADIV3       : in    std_ulogic;
          OADIV4       : in    std_ulogic;
          OAMUX0       : in    std_ulogic;
          OAMUX1       : in    std_ulogic;
          OAMUX2       : in    std_ulogic;
          DLYGLA0      : in    std_ulogic;
          DLYGLA1      : in    std_ulogic;
          DLYGLA2      : in    std_ulogic;
          DLYGLA3      : in    std_ulogic;
          DLYGLA4      : in    std_ulogic;
          OBDIV0       : in    std_ulogic;
          OBDIV1       : in    std_ulogic;
          OBDIV2       : in    std_ulogic;
          OBDIV3       : in    std_ulogic;
          OBDIV4       : in    std_ulogic;
          OBMUX0       : in    std_ulogic;
          OBMUX1       : in    std_ulogic;
          OBMUX2       : in    std_ulogic;
          DLYYB0       : in    std_ulogic;
          DLYYB1       : in    std_ulogic;
          DLYYB2       : in    std_ulogic;
          DLYYB3       : in    std_ulogic;
          DLYYB4       : in    std_ulogic;
          DLYGLB0      : in    std_ulogic;
          DLYGLB1      : in    std_ulogic;
          DLYGLB2      : in    std_ulogic;
          DLYGLB3      : in    std_ulogic;
          DLYGLB4      : in    std_ulogic;
          OCDIV0       : in    std_ulogic;
          OCDIV1       : in    std_ulogic;
          OCDIV2       : in    std_ulogic;
          OCDIV3       : in    std_ulogic;
          OCDIV4       : in    std_ulogic;
          OCMUX0       : in    std_ulogic;
          OCMUX1       : in    std_ulogic;
          OCMUX2       : in    std_ulogic;
          DLYYC0       : in    std_ulogic;
          DLYYC1       : in    std_ulogic;
          DLYYC2       : in    std_ulogic;
          DLYYC3       : in    std_ulogic;
          DLYYC4       : in    std_ulogic;
          DLYGLC0      : in    std_ulogic;
          DLYGLC1      : in    std_ulogic;
          DLYGLC2      : in    std_ulogic;
          DLYGLC3      : in    std_ulogic;
          DLYGLC4      : in    std_ulogic;
          FINDIV0      : in    std_ulogic;
          FINDIV1      : in    std_ulogic;
          FINDIV2      : in    std_ulogic;
          FINDIV3      : in    std_ulogic;
          FINDIV4      : in    std_ulogic;
          FINDIV5      : in    std_ulogic;
          FINDIV6      : in    std_ulogic;
          FBDIV0       : in    std_ulogic;
          FBDIV1       : in    std_ulogic;
          FBDIV2       : in    std_ulogic;
          FBDIV3       : in    std_ulogic;
          FBDIV4       : in    std_ulogic;
          FBDIV5       : in    std_ulogic;
          FBDIV6       : in    std_ulogic;
          FBDLY0       : in    std_ulogic;
          FBDlY1       : in    std_ulogic;
          FBDLY2       : in    std_ulogic;
          FBDLY3       : in    std_ulogic;
          FBDlY4       : in    std_ulogic;
          FBSEL0       : in    std_ulogic;
          FBSEL1       : in    std_ulogic;
          XDLYSEL      : in    std_ulogic;
          VCOSEL0      : in    std_ulogic;
          VCOSEL1      : in    std_ulogic;
          VCOSEL2      : in    std_ulogic;
          GLA          : out   std_ulogic;
          LOCK         : out   std_ulogic;
          GLB          : out   std_ulogic;
          YB           : out   std_ulogic;
          GLC          : out   std_ulogic;
          YC           : out   std_ulogic;
          SDOUT        : out   std_ulogic
        );
end component;

component DYNCCC_V2
   generic(
      VCOFREQUENCY      :  Real    := 0.0;
      f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

      TimingChecksOn    :  Boolean := True;
      InstancePath      :  STRING  := "*";
      Xon               :  Boolean := False;
      MsgOn             :  Boolean := True;

      tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKC         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SDIN         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SCLK         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SSHIFT       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SUPDATE      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_MODE         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

      tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );

      tpd_SCLK_SDOUT    : VitalDelayType01  := ( 0.100 ns, 0.100 ns );

      tsetup_SSHIFT_SCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_SSHIFT_SCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_negedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_SDIN_SCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_SDIN_SCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_negedge_posedge    : VitalDelayType := 0.000 ns;

      tpw_SUPDATE_posedge                : VitalDelayType := 0.000 ns;
      tpw_SUPDATE_negedge                : VitalDelayType := 0.000 ns;
      tpw_SCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_SCLK_negedge                   : VitalDelayType := 0.000 ns

      ); 

   port (
          CLKA         : in    std_ulogic;
          EXTFB        : in    std_ulogic;
          POWERDOWN    : in    std_ulogic;
          CLKB         : in    std_ulogic;
          CLKC         : in    std_ulogic;
          SDIN         : in    std_ulogic;
          SCLK         : in    std_ulogic;
          SSHIFT       : in    std_ulogic;
          SUPDATE      : in    std_ulogic;
          MODE         : in    std_ulogic;
          OADIV0       : in    std_ulogic;
          OADIV1       : in    std_ulogic;
          OADIV2       : in    std_ulogic;
          OADIV3       : in    std_ulogic;
          OADIV4       : in    std_ulogic;
          OAMUX0       : in    std_ulogic;
          OAMUX1       : in    std_ulogic;
          OAMUX2       : in    std_ulogic;
          DLYGLA0      : in    std_ulogic;
          DLYGLA1      : in    std_ulogic;
          DLYGLA2      : in    std_ulogic;
          DLYGLA3      : in    std_ulogic;
          DLYGLA4      : in    std_ulogic;
          OBDIV0       : in    std_ulogic;
          OBDIV1       : in    std_ulogic;
          OBDIV2       : in    std_ulogic;
          OBDIV3       : in    std_ulogic;
          OBDIV4       : in    std_ulogic;
          OBMUX0       : in    std_ulogic;
          OBMUX1       : in    std_ulogic;
          OBMUX2       : in    std_ulogic;
          DLYYB0       : in    std_ulogic;
          DLYYB1       : in    std_ulogic;
          DLYYB2       : in    std_ulogic;
          DLYYB3       : in    std_ulogic;
          DLYYB4       : in    std_ulogic;
          DLYGLB0      : in    std_ulogic;
          DLYGLB1      : in    std_ulogic;
          DLYGLB2      : in    std_ulogic;
          DLYGLB3      : in    std_ulogic;
          DLYGLB4      : in    std_ulogic;
          OCDIV0       : in    std_ulogic;
          OCDIV1       : in    std_ulogic;
          OCDIV2       : in    std_ulogic;
          OCDIV3       : in    std_ulogic;
          OCDIV4       : in    std_ulogic;
          OCMUX0       : in    std_ulogic;
          OCMUX1       : in    std_ulogic;
          OCMUX2       : in    std_ulogic;
          DLYYC0       : in    std_ulogic;
          DLYYC1       : in    std_ulogic;
          DLYYC2       : in    std_ulogic;
          DLYYC3       : in    std_ulogic;
          DLYYC4       : in    std_ulogic;
          DLYGLC0      : in    std_ulogic;
          DLYGLC1      : in    std_ulogic;
          DLYGLC2      : in    std_ulogic;
          DLYGLC3      : in    std_ulogic;
          DLYGLC4      : in    std_ulogic;
          FINDIV0      : in    std_ulogic;
          FINDIV1      : in    std_ulogic;
          FINDIV2      : in    std_ulogic;
          FINDIV3      : in    std_ulogic;
          FINDIV4      : in    std_ulogic;
          FINDIV5      : in    std_ulogic;
          FINDIV6      : in    std_ulogic;
          FBDIV0       : in    std_ulogic;
          FBDIV1       : in    std_ulogic;
          FBDIV2       : in    std_ulogic;
          FBDIV3       : in    std_ulogic;
          FBDIV4       : in    std_ulogic;
          FBDIV5       : in    std_ulogic;
          FBDIV6       : in    std_ulogic;
          FBDLY0       : in    std_ulogic;
          FBDlY1       : in    std_ulogic;
          FBDLY2       : in    std_ulogic;
          FBDLY3       : in    std_ulogic;
          FBDlY4       : in    std_ulogic;
          FBSEL0       : in    std_ulogic;
          FBSEL1       : in    std_ulogic;
          XDLYSEL      : in    std_ulogic;
          VCOSEL0      : in    std_ulogic;
          VCOSEL1      : in    std_ulogic;
          VCOSEL2      : in    std_ulogic;
          GLA          : out   std_ulogic;
          LOCK         : out   std_ulogic;
          GLB          : out   std_ulogic;
          YB           : out   std_ulogic;
          GLC          : out   std_ulogic;
          YC           : out   std_ulogic;
          SDOUT        : out   std_ulogic
        );
end component;

component SHREG
   generic(
      tipd_SDIN      : VitalDelayType01 := ( 0.0 ns, 0.0 ns );
      tipd_SCLK      : VitalDelayType01 := ( 0.0 ns, 0.0 ns );
      tipd_SSHIFT    : VitalDelayType01 := ( 0.0 ns, 0.0 ns );
      tipd_SUPDATE   : VitalDelayType01 := ( 0.0 ns, 0.0 ns );

      TimingChecksOn : Boolean := True;
      InstancePath   : STRING  := "*";
      Xon            : Boolean := False;
      MsgOn          : Boolean := True);

   port(
      SDIN           :	in    STD_ULOGIC; -- Serial data input
      SCLK           :	in    STD_ULOGIC; -- Serial Clock signal
      SSHIFT         :	in    STD_ULOGIC; -- Serial shift enable signal 
      SUPDATE        :	in    STD_ULOGIC; -- Data in SR loaded into update latch
      SDOUT          :	out   STD_ULOGIC; -- Serial data output - data from LSB of SR shifted out
      SUPDATELATCH   :  out   STD_LOGIC_VECTOR ( 80 downto 0 )); -- Configuration bits
end component;

component PLL
  generic(
     VCOFREQUENCY      :  Real    := 0.0;
     f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

     TimingChecksOn    :  Boolean          := True;
     InstancePath      :  String           := "*";
     Xon               :  Boolean          := False;
     MsgOn             :  Boolean          := True;

     tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OAMUX0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OAMUX1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OAMUX2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBMUX0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBMUX1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBMUX2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCMUX0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCMUX1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCMUX2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV5      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV6      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV5       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV6       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBSEL0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBSEL1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_XDLYSEL      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_VCOSEL0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_VCOSEL1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_VCOSEL2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );

     tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns));


  port (
     CLKA         :  in    STD_ULOGIC;
     EXTFB        :  in    STD_ULOGIC;
     POWERDOWN    :  in    STD_ULOGIC;
     OADIV0       :  in    STD_ULOGIC;
     OADIV1       :  in    STD_ULOGIC;
     OADIV2       :  in    STD_ULOGIC;
     OADIV3       :  in    STD_ULOGIC;
     OADIV4       :  in    STD_ULOGIC;
     OAMUX0       :  in    STD_ULOGIC;
     OAMUX1       :  in    STD_ULOGIC;
     OAMUX2       :  in    STD_ULOGIC;
     DLYGLA0      :  in    STD_ULOGIC;
     DLYGLA1      :  in    STD_ULOGIC;
     DLYGLA2      :  in    STD_ULOGIC;
     DLYGLA3      :  in    STD_ULOGIC;
     DLYGLA4      :  in    STD_ULOGIC;
     OBDIV0       :  in    STD_ULOGIC;
     OBDIV1       :  in    STD_ULOGIC;
     OBDIV2       :  in    STD_ULOGIC;
     OBDIV3       :  in    STD_ULOGIC;
     OBDIV4       :  in    STD_ULOGIC;
     OBMUX0       :  in    STD_ULOGIC;
     OBMUX1       :  in    STD_ULOGIC;
     OBMUX2       :  in    STD_ULOGIC;
     DLYYB0       :  in    STD_ULOGIC;
     DLYYB1       :  in    STD_ULOGIC;
     DLYYB2       :  in    STD_ULOGIC;
     DLYYB3       :  in    STD_ULOGIC;
     DLYYB4       :  in    STD_ULOGIC;
     DLYGLB0      :  in    STD_ULOGIC;
     DLYGLB1      :  in    STD_ULOGIC;
     DLYGLB2      :  in    STD_ULOGIC;
     DLYGLB3      :  in    STD_ULOGIC;
     DLYGLB4      :  in    STD_ULOGIC;
     OCDIV0       :  in    STD_ULOGIC;
     OCDIV1       :  in    STD_ULOGIC;
     OCDIV2       :  in    STD_ULOGIC;
     OCDIV3       :  in    STD_ULOGIC;
     OCDIV4       :  in    STD_ULOGIC;
     OCMUX0       :  in    STD_ULOGIC;
     OCMUX1       :  in    STD_ULOGIC;
     OCMUX2       :  in    STD_ULOGIC;
     DLYYC0       :  in    STD_ULOGIC;
     DLYYC1       :  in    STD_ULOGIC;
     DLYYC2       :  in    STD_ULOGIC;
     DLYYC3       :  in    STD_ULOGIC;
     DLYYC4       :  in    STD_ULOGIC;
     DLYGLC0      :  in    STD_ULOGIC;
     DLYGLC1      :  in    STD_ULOGIC;
     DLYGLC2      :  in    STD_ULOGIC;
     DLYGLC3      :  in    STD_ULOGIC;
     DLYGLC4      :  in    STD_ULOGIC;
     FINDIV0      :  in    STD_ULOGIC;
     FINDIV1      :  in    STD_ULOGIC;
     FINDIV2      :  in    STD_ULOGIC;
     FINDIV3      :  in    STD_ULOGIC;
     FINDIV4      :  in    STD_ULOGIC;
     FINDIV5      :  in    STD_ULOGIC;
     FINDIV6      :  in    STD_ULOGIC;
     FBDIV0       :  in    STD_ULOGIC;
     FBDIV1       :  in    STD_ULOGIC;
     FBDIV2       :  in    STD_ULOGIC;
     FBDIV3       :  in    STD_ULOGIC;
     FBDIV4       :  in    STD_ULOGIC;
     FBDIV5       :  in    STD_ULOGIC;
     FBDIV6       :  in    STD_ULOGIC;
     FBDLY0       :  in    STD_ULOGIC;
     FBDLY1       :  in    STD_ULOGIC;
     FBDLY2       :  in    STD_ULOGIC;
     FBDLY3       :  in    STD_ULOGIC;
     FBDLY4       :  in    STD_ULOGIC;
     FBSEL0       :  in    STD_ULOGIC;
     FBSEL1       :  in    STD_ULOGIC;
     XDLYSEL      :  in    STD_ULOGIC;
     VCOSEL0      :  in    STD_ULOGIC;
     VCOSEL1      :  in    STD_ULOGIC;
     VCOSEL2      :  in    STD_ULOGIC;
     GLA          :  out   STD_ULOGIC;
     LOCK         :  out   STD_ULOGIC;
     GLB          :  out   STD_ULOGIC;
     YB           :  out   STD_ULOGIC;
     GLC          :  out   STD_ULOGIC;
     YC           :  out   STD_ULOGIC);
end component;

component PLL_V2
  generic(
     VCOFREQUENCY      :  Real    := 0.0;
     f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

     TimingChecksOn    :  Boolean          := True;
     InstancePath      :  String           := "*";
     Xon               :  Boolean          := False;
     MsgOn             :  Boolean          := True;

     tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OADIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OAMUX0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OAMUX1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OAMUX2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLA4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBDIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBMUX0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBMUX1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OBMUX2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYB4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLB4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCDIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCMUX0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCMUX1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_OCMUX2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYYC4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_DLYGLC4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV3      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV4      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV5      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FINDIV6      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV5       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDIV6       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY2       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY3       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBDLY4       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBSEL0       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_FBSEL1       :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_XDLYSEL      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_VCOSEL0      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_VCOSEL1      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );
     tipd_VCOSEL2      :  VitalDelayType01 := ( 0.000 ns,0.000 ns );

     tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns);
     tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns));


  port (
     CLKA         :  in    STD_ULOGIC;
     EXTFB        :  in    STD_ULOGIC;
     POWERDOWN    :  in    STD_ULOGIC;
     OADIV0       :  in    STD_ULOGIC;
     OADIV1       :  in    STD_ULOGIC;
     OADIV2       :  in    STD_ULOGIC;
     OADIV3       :  in    STD_ULOGIC;
     OADIV4       :  in    STD_ULOGIC;
     OAMUX0       :  in    STD_ULOGIC;
     OAMUX1       :  in    STD_ULOGIC;
     OAMUX2       :  in    STD_ULOGIC;
     DLYGLA0      :  in    STD_ULOGIC;
     DLYGLA1      :  in    STD_ULOGIC;
     DLYGLA2      :  in    STD_ULOGIC;
     DLYGLA3      :  in    STD_ULOGIC;
     DLYGLA4      :  in    STD_ULOGIC;
     OBDIV0       :  in    STD_ULOGIC;
     OBDIV1       :  in    STD_ULOGIC;
     OBDIV2       :  in    STD_ULOGIC;
     OBDIV3       :  in    STD_ULOGIC;
     OBDIV4       :  in    STD_ULOGIC;
     OBMUX0       :  in    STD_ULOGIC;
     OBMUX1       :  in    STD_ULOGIC;
     OBMUX2       :  in    STD_ULOGIC;
     DLYYB0       :  in    STD_ULOGIC;
     DLYYB1       :  in    STD_ULOGIC;
     DLYYB2       :  in    STD_ULOGIC;
     DLYYB3       :  in    STD_ULOGIC;
     DLYYB4       :  in    STD_ULOGIC;
     DLYGLB0      :  in    STD_ULOGIC;
     DLYGLB1      :  in    STD_ULOGIC;
     DLYGLB2      :  in    STD_ULOGIC;
     DLYGLB3      :  in    STD_ULOGIC;
     DLYGLB4      :  in    STD_ULOGIC;
     OCDIV0       :  in    STD_ULOGIC;
     OCDIV1       :  in    STD_ULOGIC;
     OCDIV2       :  in    STD_ULOGIC;
     OCDIV3       :  in    STD_ULOGIC;
     OCDIV4       :  in    STD_ULOGIC;
     OCMUX0       :  in    STD_ULOGIC;
     OCMUX1       :  in    STD_ULOGIC;
     OCMUX2       :  in    STD_ULOGIC;
     DLYYC0       :  in    STD_ULOGIC;
     DLYYC1       :  in    STD_ULOGIC;
     DLYYC2       :  in    STD_ULOGIC;
     DLYYC3       :  in    STD_ULOGIC;
     DLYYC4       :  in    STD_ULOGIC;
     DLYGLC0      :  in    STD_ULOGIC;
     DLYGLC1      :  in    STD_ULOGIC;
     DLYGLC2      :  in    STD_ULOGIC;
     DLYGLC3      :  in    STD_ULOGIC;
     DLYGLC4      :  in    STD_ULOGIC;
     FINDIV0      :  in    STD_ULOGIC;
     FINDIV1      :  in    STD_ULOGIC;
     FINDIV2      :  in    STD_ULOGIC;
     FINDIV3      :  in    STD_ULOGIC;
     FINDIV4      :  in    STD_ULOGIC;
     FINDIV5      :  in    STD_ULOGIC;
     FINDIV6      :  in    STD_ULOGIC;
     FBDIV0       :  in    STD_ULOGIC;
     FBDIV1       :  in    STD_ULOGIC;
     FBDIV2       :  in    STD_ULOGIC;
     FBDIV3       :  in    STD_ULOGIC;
     FBDIV4       :  in    STD_ULOGIC;
     FBDIV5       :  in    STD_ULOGIC;
     FBDIV6       :  in    STD_ULOGIC;
     FBDLY0       :  in    STD_ULOGIC;
     FBDLY1       :  in    STD_ULOGIC;
     FBDLY2       :  in    STD_ULOGIC;
     FBDLY3       :  in    STD_ULOGIC;
     FBDLY4       :  in    STD_ULOGIC;
     FBSEL0       :  in    STD_ULOGIC;
     FBSEL1       :  in    STD_ULOGIC;
     XDLYSEL      :  in    STD_ULOGIC;
     VCOSEL0      :  in    STD_ULOGIC;
     VCOSEL1      :  in    STD_ULOGIC;
     VCOSEL2      :  in    STD_ULOGIC;
     GLA          :  out   STD_ULOGIC;
     LOCK         :  out   STD_ULOGIC;
     GLB          :  out   STD_ULOGIC;
     YB           :  out   STD_ULOGIC;
     GLC          :  out   STD_ULOGIC;
     YC           :  out   STD_ULOGIC);
end component;

--component CLKDIVDLY1
--     generic(
--        TimingChecksOn: Boolean := True;
--        InstancePath: STRING := "*";
--        Xon: Boolean := False;
--        MsgOn: Boolean := True;
--        tipd_CLK         :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns );
--        tpd_CLK_Y         :  VitalDelayType01 := (  0.1 ns,0.1 ns ));
--
--
--     port (
--        CLK         : in    STD_ULOGIC;
--        ODIV0       : in    STD_ULOGIC;
--        ODIV1       : in    STD_ULOGIC;
--        ODIV2       : in    STD_ULOGIC;
--        ODIV3       : in    STD_ULOGIC;
--        ODIV4       : in    STD_ULOGIC;
--        DLYY0       : in    STD_ULOGIC;
--        DLYY1       : in    STD_ULOGIC;
--        DLYY2       : in    STD_ULOGIC;
--        DLYY3       : in    STD_ULOGIC;
--        DLYY4       : in    STD_ULOGIC;
--        DLYGL0       : in    STD_ULOGIC;
--        DLYGL1       : in    STD_ULOGIC;
--        DLYGL2       : in    STD_ULOGIC;
--        DLYGL3       : in    STD_ULOGIC;
--        DLYGL4       : in    STD_ULOGIC;
--        GL           : out   STD_ULOGIC;
--        Y            : out   STD_ULOGIC);
-- 
--end component;

--component CLKDIVDLY
--     generic(
--        TimingChecksOn: Boolean := True;
--        InstancePath: STRING := "*";
--        Xon: Boolean := False;
--        MsgOn: Boolean := True;
--        tipd_CLK         :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns ));
--
--     port (
--        CLK         : in    STD_ULOGIC;
--        ODIV0       : in    STD_ULOGIC;
--        ODIV1       : in    STD_ULOGIC;
--        ODIV2       : in    STD_ULOGIC;
--        ODIV3       : in    STD_ULOGIC;
--        ODIV4       : in    STD_ULOGIC;
--        DLYGL0       : in    STD_ULOGIC;
--        DLYGL1       : in    STD_ULOGIC;
--        DLYGL2       : in    STD_ULOGIC;
--        DLYGL3       : in    STD_ULOGIC;
--        DLYGL4       : in    STD_ULOGIC;
--        GL           : out   STD_ULOGIC
--          );
--
--end component;

component CLKDLY
    generic(
        TimingChecksOn: Boolean := True;
        InstancePath: STRING := "*";
        Xon: Boolean := False;
        MsgOn: Boolean := True;
        tipd_CLK          :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns )
        );

     port (
        CLK          : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL           : out   STD_ULOGIC
          );

end component;

component CLKDLYIO
    generic(
        TimingChecksOn    : Boolean := True;
        InstancePath      : STRING  := "*";
        Xon               : Boolean := False;
        MsgOn             : Boolean := True;
        tipd_CLK          : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL0       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL1       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL2       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL3       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL4       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tpd_CLK_GL        : VitalDelayType01  := (  0.1 ns,0.1 ns )
        ); 
    port (
        CLK          : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL           : out   STD_ULOGIC
        );
end component;

component CLKDLYINT
    generic(
        TimingChecksOn    : Boolean := True;
        InstancePath      : STRING  := "*";
        Xon               : Boolean := False;
        MsgOn             : Boolean := True;
        tipd_CLK          : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL0       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL1       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL2       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL3       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tipd_DLYGL4       : VitalDelayType01  := (  0.0 ns,0.0 ns );
        tpd_CLK_GL        : VitalDelayType01  := (  0.1 ns,0.1 ns )
        );
    port (
        CLK          : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL           : out   STD_ULOGIC
        );
end component;

component RAM4K9
   generic (
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;
      MEMORYFILE       : String  := "";
      WARNING_MSGS_ON  : Boolean := True;
           
      tipd_ADDRA11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA8       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA7       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA6       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA5       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA4       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA3       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA2       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB8       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB7       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB6       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB5       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB4       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB3       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB2       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHA1     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHA0     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHB1     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHB0     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PIPEA       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PIPEB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WMODEA      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WMODEB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_BLKA        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_BLKB        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WENA        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WENB        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLKA        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLKB        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RESET       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLKA_DOUTA8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA8 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA7 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA6 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA5 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA4 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA3 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA2 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA1 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA0 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB8 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB7 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB6 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB5 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB4 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB3 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB2 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB1 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB0 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tsetup_DINA8_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA8_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA7_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA7_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA6_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA6_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA5_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA5_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA4_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA4_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA3_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA3_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA2_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA2_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA1_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA1_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA0_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINA0_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB8_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB8_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB7_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB7_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB6_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB6_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB5_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB5_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB4_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB4_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB3_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB3_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB2_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB2_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB1_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB1_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB0_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_DINB0_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA8_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA8_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA7_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA7_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA6_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA6_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA5_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA5_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA4_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA4_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA3_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA3_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA2_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA2_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA1_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA1_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA0_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINA0_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB8_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB8_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB7_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB7_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB6_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB6_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB5_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB5_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB4_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB4_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB3_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB3_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB2_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB2_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB1_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB1_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB0_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DINB0_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_ADDRA11_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA11_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA10_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA10_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA9_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA9_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA8_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA8_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA7_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA7_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA6_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA6_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA5_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA5_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA4_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA4_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA3_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA3_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA2_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA2_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA1_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA1_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA0_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRA0_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA11_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA11_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA10_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA10_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA9_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA9_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA8_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA8_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA7_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA7_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA6_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA6_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA5_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA5_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA4_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA4_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA3_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA3_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA2_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA2_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA1_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA1_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA0_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRA0_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_ADDRB11_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB11_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB10_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB10_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB9_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB9_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB8_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB8_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB7_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB7_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB6_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB6_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB5_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB5_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB4_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB4_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB3_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB3_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB2_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB2_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB1_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB1_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB0_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB0_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB11_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB11_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB10_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB10_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB9_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB9_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB8_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB8_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB7_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB7_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB6_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB6_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB5_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB5_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB4_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB4_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB3_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB3_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB2_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB2_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB1_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB1_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB0_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_ADDRB0_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WENA_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WENA_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_BLKA_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_BLKA_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WMODEA_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WMODEA_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_PIPEA_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_PIPEA_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_WENA_CLKA_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WENA_CLKA_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_BLKA_CLKA_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_BLKA_CLKA_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WMODEA_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_WMODEA_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_PIPEA_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_PIPEA_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WENB_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WENB_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_BLKB_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_BLKB_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WMODEB_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WMODEB_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_PIPEB_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_PIPEB_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB1_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB1_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHB1_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WIDTHB1_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB0_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB0_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHB0_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WIDTHB0_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;

      tsetup_WIDTHA1_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WIDTHA1_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHA1_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WIDTHA1_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WIDTHA0_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WIDTHA0_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHA0_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WIDTHA0_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;

      thold_WENB_CLKB_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WENB_CLKB_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_BLKB_CLKB_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_BLKB_CLKB_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WMODEB_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_WMODEB_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_PIPEB_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_PIPEB_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      
      tpw_CLKA_posedge                     : VitalDelayType := 0.000 ns;
      tpw_CLKA_negedge                     : VitalDelayType := 0.000 ns;
      tpw_CLKB_posedge                     : VitalDelayType := 0.000 ns;
      tpw_CLKB_negedge                     : VitalDelayType := 0.000 ns;
      trecovery_RESET_CLKA_posedge_posedge : VitalDelayType := 0.000 ns;
      trecovery_RESET_CLKB_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_RESET_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RESET_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      tpw_RESET_negedge                    : VitalDelayType := 0.000 ns
     );

   port (
      ADDRA11       : IN STD_ULOGIC ;
      ADDRA10       : IN STD_ULOGIC ;
      ADDRA9        : IN STD_ULOGIC ;
      ADDRA8        : IN STD_ULOGIC ;
      ADDRA7        : IN STD_ULOGIC ;
      ADDRA6        : IN STD_ULOGIC ;
      ADDRA5        : IN STD_ULOGIC ;
      ADDRA4        : IN STD_ULOGIC ;
      ADDRA3        : IN STD_ULOGIC ;
      ADDRA2        : IN STD_ULOGIC ;
      ADDRA1        : IN STD_ULOGIC ;
      ADDRA0        : IN STD_ULOGIC ;
      ADDRB11       : IN STD_ULOGIC ;
      ADDRB10       : IN STD_ULOGIC ;
      ADDRB9        : IN STD_ULOGIC ;
      ADDRB8        : IN STD_ULOGIC ;
      ADDRB7        : IN STD_ULOGIC ;
      ADDRB6        : IN STD_ULOGIC ;
      ADDRB5        : IN STD_ULOGIC ;
      ADDRB4        : IN STD_ULOGIC ;
      ADDRB3        : IN STD_ULOGIC ;
      ADDRB2        : IN STD_ULOGIC ;
      ADDRB1        : IN STD_ULOGIC ;
      ADDRB0        : IN STD_ULOGIC ;
      DINA8         : IN STD_ULOGIC ;
      DINA7         : IN STD_ULOGIC ;
      DINA6         : IN STD_ULOGIC ;
      DINA5         : IN STD_ULOGIC ;
      DINA4         : IN STD_ULOGIC ;
      DINA3         : IN STD_ULOGIC ;
      DINA2         : IN STD_ULOGIC ;
      DINA1         : IN STD_ULOGIC ;
      DINA0         : IN STD_ULOGIC ; 
      DINB8         : IN STD_ULOGIC ;
      DINB7         : IN STD_ULOGIC ;
      DINB6         : IN STD_ULOGIC ;
      DINB5         : IN STD_ULOGIC ;
      DINB4         : IN STD_ULOGIC ;
      DINB3         : IN STD_ULOGIC ;
      DINB2         : IN STD_ULOGIC ;
      DINB1         : IN STD_ULOGIC ;
      DINB0         : IN STD_ULOGIC ;
      WIDTHA1       : IN STD_ULOGIC ;
      WIDTHA0       : IN STD_ULOGIC ;
      WIDTHB1       : IN STD_ULOGIC ;
      WIDTHB0       : IN STD_ULOGIC ;
      PIPEA         : IN STD_ULOGIC ;
      PIPEB         : IN STD_ULOGIC ;
      WMODEA        : IN STD_ULOGIC ;
      WMODEB        : IN STD_ULOGIC ;
      BLKA          : IN STD_ULOGIC ;
      BLKB          : IN STD_ULOGIC ;
      WENA          : IN STD_ULOGIC ;
      WENB          : IN STD_ULOGIC ;
      CLKA          : IN STD_ULOGIC ;
      CLKB          : IN STD_ULOGIC ;
      RESET         : IN STD_ULOGIC ;
      DOUTA8        : OUT STD_ULOGIC ;
      DOUTA7        : OUT STD_ULOGIC ;
      DOUTA6        : OUT STD_ULOGIC ;
      DOUTA5        : OUT STD_ULOGIC ;
      DOUTA4        : OUT STD_ULOGIC ;
      DOUTA3        : OUT STD_ULOGIC ;
      DOUTA2        : OUT STD_ULOGIC ;
      DOUTA1        : OUT STD_ULOGIC ;
      DOUTA0        : OUT STD_ULOGIC ;
      DOUTB8        : OUT STD_ULOGIC ;
      DOUTB7        : OUT STD_ULOGIC ;
      DOUTB6        : OUT STD_ULOGIC ;
      DOUTB5        : OUT STD_ULOGIC ;
      DOUTB4        : OUT STD_ULOGIC ;
      DOUTB3        : OUT STD_ULOGIC ;
      DOUTB2        : OUT STD_ULOGIC ;
      DOUTB1        : OUT STD_ULOGIC ;
      DOUTB0        : OUT STD_ULOGIC
     );

end component;


component RAM512X18
   generic (
      TimingChecksOn  : Boolean := True;
      InstancePath    : String  := "*";
      Xon             : Boolean := False;
      MsgOn           : Boolean := True;
      MEMORYFILE      : String  := "";
      WARNING_MSGS_ON : Boolean := True;

      tipd_RADDR8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD17      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD16      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD15      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD14      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD13      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD12      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD11      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD10      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD9       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD8       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD7       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD6       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD5       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD4       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD3       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD2       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WEN       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WCLK      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REN       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RCLK      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PIPE      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RESET     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      
      tpd_RCLK_RD17  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RCLK_RD16  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD15  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD14  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD13  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD12  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD11  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD10  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD9   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD8   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD7   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD6   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD5   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD4   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD3   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD2   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD1   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD0   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      
      tsetup_WD17_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD17_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD16_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD16_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD15_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD15_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD14_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD14_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD13_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD13_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD12_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD12_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD11_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD11_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD10_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD10_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD9_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD9_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD8_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD8_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD7_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD7_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD6_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD6_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD5_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD5_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD4_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD4_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD17_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD17_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD16_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD16_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WADDR8_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR8_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR7_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR7_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR6_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR6_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR5_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR5_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR4_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR4_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR3_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR3_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR2_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR2_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR1_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR1_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR0_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR0_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_WADDR8_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;    
      thold_WADDR8_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR7_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR7_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR6_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR6_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR5_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR5_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR4_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR4_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WW1_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WW1_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WW0_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WW0_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WEN_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WEN_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_WW1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WW1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WW0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WW0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WEN_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WEN_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_RADDR8_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;    
      tsetup_RADDR8_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR7_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR7_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR6_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR6_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR5_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR5_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR4_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR4_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR3_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR3_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR2_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR2_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR1_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR1_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR0_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR0_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_RADDR8_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;    
      thold_RADDR8_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR7_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR7_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR6_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR6_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR5_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR5_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR4_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR4_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR3_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR3_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR2_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR2_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR1_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR1_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR0_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR0_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_RW1_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_RW1_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_RW0_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_RW0_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_REN_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_REN_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_RW1_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RW1_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RW0_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RW0_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_REN_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_REN_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;      
      tsetup_PIPE_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_PIPE_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_PIPE_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_PIPE_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tpw_WCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_WCLK_negedge                   : VitalDelayType := 0.000 ns;
      tpw_RCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_RCLK_negedge                   : VitalDelayType := 0.000 ns;
      trecovery_RESET_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      trecovery_RESET_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_RESET_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RESET_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tpw_RESET_negedge                    : VitalDelayType := 0.000 ns
     );

     port (
           RADDR8        : IN STD_ULOGIC ;
           RADDR7        : IN STD_ULOGIC ;
           RADDR6        : IN STD_ULOGIC ;
           RADDR5        : IN STD_ULOGIC ;
           RADDR4        : IN STD_ULOGIC ;
           RADDR3        : IN STD_ULOGIC ;
           RADDR2        : IN STD_ULOGIC ;
           RADDR1        : IN STD_ULOGIC ;  
           RADDR0        : IN STD_ULOGIC ;
           WADDR8        : IN STD_ULOGIC ;
           WADDR7        : IN STD_ULOGIC ;
           WADDR6        : IN STD_ULOGIC ;
           WADDR5        : IN STD_ULOGIC ;
           WADDR4        : IN STD_ULOGIC ;
           WADDR3        : IN STD_ULOGIC ;
           WADDR2        : IN STD_ULOGIC ;
           WADDR1        : IN STD_ULOGIC ;
           WADDR0        : IN STD_ULOGIC ;
           WD17          : IN STD_ULOGIC ;
           WD16          : IN STD_ULOGIC ;
           WD15          : IN STD_ULOGIC ;
           WD14          : IN STD_ULOGIC ;
           WD13          : IN STD_ULOGIC ;
           WD12          : IN STD_ULOGIC ;
           WD11          : IN STD_ULOGIC ;
           WD10          : IN STD_ULOGIC ;
           WD9           : IN STD_ULOGIC ;
           WD8           : IN STD_ULOGIC ;
           WD7           : IN STD_ULOGIC ;
           WD6           : IN STD_ULOGIC ;
           WD5           : IN STD_ULOGIC ;
           WD4           : IN STD_ULOGIC ;
           WD3           : IN STD_ULOGIC ;
           WD2           : IN STD_ULOGIC ;
           WD1           : IN STD_ULOGIC ;
           WD0           : IN STD_ULOGIC ;
           WW1           : IN STD_ULOGIC ;
           WW0           : IN STD_ULOGIC ;
           WEN           : IN STD_ULOGIC ;
           WCLK          : IN STD_ULOGIC ;
           RW1           : IN STD_ULOGIC ;
           RW0           : IN STD_ULOGIC ;
           REN           : IN STD_ULOGIC ;
           RCLK          : IN STD_ULOGIC ;
           PIPE          : IN STD_ULOGIC ;
           RESET         : IN STD_ULOGIC ;
           RD17          : OUT STD_ULOGIC ;
           RD16          : OUT STD_ULOGIC ;
           RD15          : OUT STD_ULOGIC ;
           RD14          : OUT STD_ULOGIC ;
           RD13          : OUT STD_ULOGIC ;
           RD12          : OUT STD_ULOGIC ;
           RD11          : OUT STD_ULOGIC ;
           RD10          : OUT STD_ULOGIC ;
           RD9           : OUT STD_ULOGIC ;
           RD8           : OUT STD_ULOGIC ;
           RD7           : OUT STD_ULOGIC ;
           RD6           : OUT STD_ULOGIC ;
           RD5           : OUT STD_ULOGIC ;
           RD4           : OUT STD_ULOGIC ;
           RD3           : OUT STD_ULOGIC ;
           RD2           : OUT STD_ULOGIC ;
           RD1           : OUT STD_ULOGIC ;
           RD0           : OUT STD_ULOGIC
  );

end component;

component FIFO4K18 
  generic(
          TimingChecksOn : Boolean := True;
          InstancePath   : String  := "*";
          Xon            : Boolean := False;
          MsgOn          : Boolean := True;

          tipd_AEVAL11  : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL10  : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL9   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL8   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL7   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL6   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL5   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL4   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AEVAL0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL11  : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL10  : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL9   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL8   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL7   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL6   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL5   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL4   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL3   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL2   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL1   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_AFVAL0   : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_REN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RBLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WEN      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WBLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WCLK     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RESET    : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RPIPE    : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_RW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WW2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WW1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WW0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_ESTOP    : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_FSTOP    : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD17     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD16     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD15     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD14     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD13     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD12     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tipd_WD0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
          tpd_RCLK_RD17     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD16     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD15     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD14     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD13     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD12     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD11     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD10     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD9      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD8      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD7      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD6      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD5      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD4      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD3      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD2      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD1      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_RD0      : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RCLK_EMPTY    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
          tpd_RCLK_AEMPTY   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
          tpd_RCLK_AFULL    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
          tpd_WCLK_FULL     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
          tpd_WCLK_AFULL    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
          tpd_WCLK_AEMPTY   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
          tpd_RESET_RD17    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD16    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD15    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD14    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD13    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD12    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD11    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD10    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD9     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD8     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD7     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD6     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD5     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD4     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD3     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD2     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD1     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_RD0     : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_EMPTY   : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_AEMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_FULL    : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tpd_RESET_AFULL   : VitalDelayType01 := (0.100 ns, 0.100 ns);
          tsetup_WD17_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD17_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD16_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD16_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD15_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD15_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD14_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD14_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD13_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD13_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD12_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD12_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD11_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD11_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD10_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD10_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD9_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD9_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD8_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD8_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD7_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD7_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD6_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD6_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD5_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD5_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD4_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD4_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD3_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD3_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD2_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD2_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD1_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD1_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD0_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WD0_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD17_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD17_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD16_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD16_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD15_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD15_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD14_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD14_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD13_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD13_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD12_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD12_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD11_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD11_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD10_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD10_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD9_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD9_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD8_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD8_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD7_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD7_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD6_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD6_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD5_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD5_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD4_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD4_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD3_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD3_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD2_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD2_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD1_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD1_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD0_WCLK_posedge_posedge              : VitalDelayType := 0.000 ns;
          thold_WD0_WCLK_negedge_posedge              : VitalDelayType := 0.000 ns;
          tsetup_WEN_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WEN_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WBLK_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WBLK_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WEN_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WEN_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WBLK_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WBLK_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_REN_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_REN_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RBLK_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RBLK_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_REN_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_REN_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RBLK_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RBLK_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_FSTOP_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_FSTOP_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_ESTOP_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_ESTOP_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_FSTOP_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_FSTOP_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_ESTOP_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_ESTOP_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WW2_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WW2_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WW1_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WW1_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WW0_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_WW0_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WW2_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WW2_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WW1_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WW1_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WW0_WCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_WW0_WCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RW2_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RW2_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RW1_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RW1_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RW0_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          tsetup_RW0_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RW2_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RW2_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RW1_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RW1_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RW0_RCLK_posedge_posedge             : VitalDelayType := 0.000 ns;
          thold_RW0_RCLK_negedge_posedge             : VitalDelayType := 0.000 ns;
          tpw_WCLK_posedge                           : VitalDelayType := 0.000 ns;
          tpw_WCLK_negedge                           : VitalDelayType := 0.000 ns;
          tperiod_WCLK                               : VitalDelayType := 0.000 ns;                                   
          tpw_RCLK_posedge                           : VitalDelayType := 0.000 ns;
          tpw_RCLK_negedge                           : VitalDelayType := 0.000 ns;
          tperiod_RCLK                               : VitalDelayType := 0.000 ns;                                   
          trecovery_RESET_RCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
          trecovery_RESET_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
          thold_RESET_RCLK_posedge_posedge           : VitalDelayType := 0.000 ns;
          thold_RESET_WCLK_posedge_posedge           : VitalDelayType := 0.000 ns;
          tpw_RESET_negedge                          : VitalDelayType := 0.000 ns

         );

port (
          AEVAL11       : IN STD_ULOGIC ;
          AEVAL10       : IN STD_ULOGIC ;
          AEVAL9       : IN STD_ULOGIC ;
          AEVAL8       : IN STD_ULOGIC ;
          AEVAL7       : IN STD_ULOGIC ;
          AEVAL6       : IN STD_ULOGIC ;
          AEVAL5       : IN STD_ULOGIC ;
          AEVAL4       : IN STD_ULOGIC ;
          AEVAL3       : IN STD_ULOGIC ;
          AEVAL2       : IN STD_ULOGIC ;
          AEVAL1       : IN STD_ULOGIC ;
          AEVAL0       : IN STD_ULOGIC ;
          AFVAL11       : IN STD_ULOGIC ;
          AFVAL10       : IN STD_ULOGIC ;
          AFVAL9       : IN STD_ULOGIC ;
          AFVAL8       : IN STD_ULOGIC ;
          AFVAL7       : IN STD_ULOGIC ;
          AFVAL6       : IN STD_ULOGIC ;
          AFVAL5       : IN STD_ULOGIC ;
          AFVAL4       : IN STD_ULOGIC ;
          AFVAL3       : IN STD_ULOGIC ;
          AFVAL2       : IN STD_ULOGIC ;
          AFVAL1       : IN STD_ULOGIC ;
          AFVAL0       : IN STD_ULOGIC ;
          REN          : IN STD_ULOGIC ;
          RBLK          : IN STD_ULOGIC ;
          RCLK          : IN STD_ULOGIC ;
          RESET         : IN STD_ULOGIC ;
          RPIPE         : IN STD_ULOGIC ;
          WEN           : IN STD_ULOGIC ;
          WBLK          : IN STD_ULOGIC ;
          WCLK          : IN STD_ULOGIC ;
          RW2           : IN STD_ULOGIC ;
          RW1           : IN STD_ULOGIC ;
          RW0           : IN STD_ULOGIC ;
          WW2           : IN STD_ULOGIC ;
          WW1           : IN STD_ULOGIC ;
          WW0           : IN STD_ULOGIC ;
          ESTOP         : IN STD_ULOGIC ;
          FSTOP         : IN STD_ULOGIC ;
          WD17          : IN STD_ULOGIC ;
          WD16          : IN STD_ULOGIC ;
          WD15          : IN STD_ULOGIC ;
          WD14          : IN STD_ULOGIC ;
          WD13          : IN STD_ULOGIC ;
          WD12          : IN STD_ULOGIC ;
          WD11          : IN STD_ULOGIC ;
          WD10          : IN STD_ULOGIC ;
          WD9           : IN STD_ULOGIC ;
          WD8           : IN STD_ULOGIC ;
          WD7           : IN STD_ULOGIC ;
          WD6           : IN STD_ULOGIC ;
          WD5           : IN STD_ULOGIC ;
          WD4           : IN STD_ULOGIC ;
          WD3           : IN STD_ULOGIC ;
          WD2           : IN STD_ULOGIC ;
          WD1           : IN STD_ULOGIC ;
          WD0           : IN STD_ULOGIC ;
          RD17          : OUT STD_ULOGIC ;
          RD16          : OUT STD_ULOGIC ;
          RD15          : OUT STD_ULOGIC ;
          RD14          : OUT STD_ULOGIC ;
          RD13          : OUT STD_ULOGIC ;
          RD12          : OUT STD_ULOGIC ;
          RD11          : OUT STD_ULOGIC ;
          RD10          : OUT STD_ULOGIC ;
          RD9           : OUT STD_ULOGIC ;
          RD8           : OUT STD_ULOGIC ;
          RD7           : OUT STD_ULOGIC ;
          RD6           : OUT STD_ULOGIC ;
          RD5           : OUT STD_ULOGIC ;
          RD4           : OUT STD_ULOGIC ;
          RD3           : OUT STD_ULOGIC ;
          RD2           : OUT STD_ULOGIC ;
          RD1           : OUT STD_ULOGIC ;
          RD0           : OUT STD_ULOGIC ;
          FULL          : OUT STD_ULOGIC ;
          AFULL         : OUT STD_ULOGIC ;
          EMPTY         : OUT STD_ULOGIC ;
          AEMPTY        : OUT STD_ULOGIC
         );


end component;


 
component DDR_OUT 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_Q      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLK_Q     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tsetup_DR_CLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_CLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                thold_CLR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_CLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                CLK            :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                Q               :  out    STD_ULOGIC);
 end component;

  component DDR_REG 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_QR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_QF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLK_QR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLK_QF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tsetup_D_CLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_D_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_D_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_D_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_CLR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_CLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_D        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                CLK            :   in    STD_ULOGIC;
                D             :  in    STD_ULOGIC;
                QF               :  out    STD_ULOGIC;
                QR               :  out    STD_ULOGIC);

 end component;

------ Component IOBI_ID_OB_EB ------
 component IOBI_ID_OB_EB
   generic (
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;

      tipd_D           : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E           : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ICLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_YIN         : VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_D_DOUT       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_E_EOUT       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLR_YR       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLR_YF       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_ICLK_YR      : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_ICLK_YF      : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_YIN_ICLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_YIN_ICLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_negedge_posedge     : VitalDelayType := 0.000 ns;

      tsetup_YIN_ICLK_posedge_negedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_posedge_negedge     : VitalDelayType := 0.000 ns;
      tsetup_YIN_ICLK_negedge_negedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_negedge_negedge     : VitalDelayType := 0.000 ns;

      trecovery_CLR_ICLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_CLR_ICLK_negedge_posedge     : VitalDelayType := 0.000 ns;

      tpw_ICLK_posedge                   :  VitalDelayType := 0.000 ns;
      tpw_ICLK_negedge                   :  VitalDelayType := 0.000 ns;
      tperiod_ICLK_posedge               :  VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                    :  VitalDelayType := 0.000 ns
     );


   port (
      D             :  in    std_ulogic;
      CLR           :  in    std_ulogic;
      E             :  in    std_ulogic;
      ICLK          :  in    std_ulogic;
      YIN           :  in    std_ulogic;
      DOUT          :  out   std_ulogic;
      EOUT          :  out   std_ulogic;
      YR            :  out   std_ulogic;
      YF            :  out   std_ulogic
     );
 end component;

 component IOBI_ID_OD_EB 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_EOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_YIN_ICLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_YIN_ICLK_posedge_negedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;



                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                thold_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_ICLK_posedge    :  VitalDelayType := 0.000 ns;

                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;

                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_YIN        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_ICLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                ICLK            :   in    STD_ULOGIC;
                YIN             :   in    STD_ULOGIC;
                E               :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                YR               :  out    STD_ULOGIC;
                YF               :  out    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 end component;

 component IOBI_ID_OD_ERC 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_EOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_EOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tpd_CLR_YR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_YIN_ICLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_YIN_ICLK_posedge_negedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_E_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
    
                
                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                thold_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_ICLK_posedge    :  VitalDelayType := 0.000 ns;

                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge    :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_YIN        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_ICLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                ICLK            :   in    STD_ULOGIC;
                YIN             :   in    STD_ULOGIC;
                E               :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                YR               :  out    STD_ULOGIC;
                YF               :  out    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 end component;


 component IOIN_ID 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_YR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_YIN_ICLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_posedge_negedge  :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_negedge  :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;

                thold_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_ICLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_YIN        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_ICLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));

 
  port(
                CLR             :   in    STD_ULOGIC;
                ICLK            :   in    STD_ULOGIC;
                YIN             :  in    STD_ULOGIC;
                YF               :  out    STD_ULOGIC;
                YR               :  out    STD_ULOGIC);

 end component;


 component IOTRI_OD_EB 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_EOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));




  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                E              :  in    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 end component;

 component IOTRI_OD_ERC 
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_EOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_EOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_E_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;


                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                E             :  in    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 end component;

------ Component AND2 ------
 component AND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND2A ------
 component AND2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND2B ------
 component AND2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND2FT ------
 component AND2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3 ------
 component AND3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3A ------
 component AND3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3B ------
 component AND3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3C ------
 component AND3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO12 ------
 component AO12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO13 ------
 component AO13
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO14 ------
 component AO14
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO15 ------
 component AO15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO16 ------
 component AO16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO17 ------
 component AO17
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO18 ------
 component AO18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1 ------
 component AO1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1A ------
 component AO1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1B ------
 component AO1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1C ------
 component AO1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1D ------
 component AO1D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO1E ------
 component AO1E
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1 ------
 component AOI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1A ------
 component AOI1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1B ------
 component AOI1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1C ------
 component AOI1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI1D ------
 component AOI1D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI5 ------
 component AOI5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1 ------
 component AX1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1A ------
 component AX1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1B ------
 component AX1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1C ------
 component AX1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1D ------
 component AX1D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AX1E ------
 component AX1E
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO1 ------
 component AXO1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO2 ------
 component AXO2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO3 ------
 component AXO3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO5 ------
 component AXO5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO6 ------
 component AXO6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXO7 ------
 component AXO7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI1 ------
 component AXOI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI2 ------
 component AXOI2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI3 ------
 component AXOI3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI4 ------
 component AXOI4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI5 ------
 component AXOI5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AXOI7 ------
 component AXOI7
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF ------
 component BIBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_12 ------
 component BIBUF_F_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_12D ------
 component BIBUF_F_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_12U ------
 component BIBUF_F_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_16 ------
 component BIBUF_F_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_16D ------
 component BIBUF_F_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_16U ------
 component BIBUF_F_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_8 ------
 component BIBUF_F_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_8D ------
 component BIBUF_F_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_8U ------
 component BIBUF_F_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_24 ------
 component BIBUF_F_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_24D ------
 component BIBUF_F_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_24U ------
 component BIBUF_F_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS15 ------
 component BIBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS15D ------
 component BIBUF_LVCMOS15D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS15U ------
 component BIBUF_LVCMOS15U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component BIBUF_LVCMOS12 ------
 component BIBUF_LVCMOS12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS12D ------
 component BIBUF_LVCMOS12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS12U ------
 component BIBUF_LVCMOS12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS18 ------
 component BIBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS18D ------
 component BIBUF_LVCMOS18D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS18U ------
 component BIBUF_LVCMOS18U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS25 ------
 component BIBUF_LVCMOS25
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS25D ------
 component BIBUF_LVCMOS25D
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS33 ------
 component BIBUF_LVCMOS33
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS25U ------
 component BIBUF_LVCMOS25U
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS33D ------
 component BIBUF_LVCMOS33D
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS33U ------
 component BIBUF_LVCMOS33U
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS5 ------
 component BIBUF_LVCMOS5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS5D ------
 component BIBUF_LVCMOS5D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_LVCMOS5U ------
 component BIBUF_LVCMOS5U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


component BIBUF_LVDS
    generic(
       TimingChecksOn : Boolean  := True;
       Xon            : Boolean  := False;
       InstancePath   : STRING   := "*";
       MsgOn          : Boolean  := True;

                tpw_D_posedge    : VitalDelayType    := 0.000 ns;
                tpw_D_negedge    : VitalDelayType    := 0.000 ns;
                tpw_E_posedge    : VitalDelayType    := 0.000 ns;
                tpw_E_negedge    : VitalDelayType    := 0.000 ns;
                tpw_PADP_negedge : VitalDelayType    := 0.000 ns;
                tpw_PADP_posedge : VitalDelayType    := 0.000 ns;
                tpw_PADN_negedge : VitalDelayType    := 0.000 ns;
                tpw_PADN_posedge : VitalDelayType    := 0.000 ns;

                tpd_D_PADP       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADP       : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_D_PADN       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADN       : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_PADP_Y       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_PADN_Y       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_D_Y          : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_Y          : VitalDelayType01  := (0.100 ns, 0.100 ns);

                tipd_D           : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_E           : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PADP        : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PADN        : VitalDelayType01  := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PADP            : inout STD_ULOGIC;
                PADN            : inout STD_ULOGIC;
                Y               : out   STD_ULOGIC);
end component;


------ Component BIBUF_PCI ------
 component BIBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_PCIX ------
 component BIBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_12 ------
 component BIBUF_S_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_12D ------
 component BIBUF_S_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_12U ------
 component BIBUF_S_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_16 ------
 component BIBUF_S_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_16D ------
 component BIBUF_S_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_16U ------
 component BIBUF_S_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_8 ------
 component BIBUF_S_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_8D ------
 component BIBUF_S_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_8U ------
 component BIBUF_S_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_24 ------
 component BIBUF_S_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_24D ------
 component BIBUF_S_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_24U ------
 component BIBUF_S_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF ------
 component CLKBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS15 ------
 component CLKBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component CLKBUF_LVCMOS12 ------
 component CLKBUF_LVCMOS12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS18 ------
 component CLKBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS25 ------
 component CLKBUF_LVCMOS25
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS33 ------
 component CLKBUF_LVCMOS33
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVCMOS5 ------
 component CLKBUF_LVCMOS5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_LVDS ------
  


component CLKBUF_LVDS
     generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
 end component;

------ Component CLKBUF_LVPECL ------
 component CLKBUF_LVPECL
     generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

 end component;

------ Component CLKBUF_PCI ------
 component CLKBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBUF_PCIX ------
 component CLKBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component DFI0 ------
 component DFI0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0C0 ------
 component DFI0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0C1 ------
 component DFI0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E0 ------
 component DFI0E0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E0C0 ------
 component DFI0E0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E0C1 ------
 component DFI0E0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E0P0 ------
 component DFI0E0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E0P1 ------
 component DFI0E0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E1 ------
 component DFI0E1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E1C0 ------
 component DFI0E1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E1C1 ------
 component DFI0E1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E1P0 ------
 component DFI0E1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0E1P1 ------
 component DFI0E1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0P0 ------
 component DFI0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0P1 ------
 component DFI0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI0P1C1 ------
 component DFI0P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1 ------
 component DFI1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1C0 ------
 component DFI1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1C1 ------
 component DFI1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E0 ------
 component DFI1E0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E0C0 ------
 component DFI1E0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E0C1 ------
 component DFI1E0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E0P0 ------
 component DFI1E0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E0P1 ------
 component DFI1E0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E1 ------
 component DFI1E1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E1C0 ------
 component DFI1E1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E1C1 ------
 component DFI1E1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E1P0 ------
 component DFI1E1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1E1P1 ------
 component DFI1E1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1P0 ------
 component DFI1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1P1 ------
 component DFI1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFI1P1C1 ------
 component DFI1P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DFN0 ------
 component DFN0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0C0 ------
 component DFN0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0C1 ------
 component DFN0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E0 ------
 component DFN0E0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E0C0 ------
 component DFN0E0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E0C1 ------
 component DFN0E0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E0P0 ------
 component DFN0E0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E0P1 ------
 component DFN0E0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E1 ------
 component DFN0E1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E1C0 ------
 component DFN0E1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E1C1 ------
 component DFN0E1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E1P0 ------
 component DFN0E1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0E1P1 ------
 component DFN0E1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0P0 ------
 component DFN0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0P1 ------
 component DFN0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN0P1C1 ------
 component DFN0P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1 ------
 component DFN1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1C0 ------
 component DFN1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1C1 ------
 component DFN1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E0 ------
 component DFN1E0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E0C0 ------
 component DFN1E0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E0C1 ------
 component DFN1E0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E0P0 ------
 component DFN1E0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E0P1 ------
 component DFN1E0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E1 ------
 component DFN1E1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E1C0 ------
 component DFN1E1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E1C1 ------
 component DFN1E1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E1P0 ------
 component DFN1E1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1E1P1 ------
 component DFN1E1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1P0 ------
 component DFN1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1P1 ------
 component DFN1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFN1P1C1 ------
 component DFN1P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLI0 ------
 component DLI0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI0C0 ------
 component DLI0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI0C1 ------
 component DLI0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI0P0 ------
 component DLI0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI0P1 ------
 component DLI0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI0P1C1 ------
 component DLI0P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI1 ------
 component DLI1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI1C0 ------
 component DLI1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI1C1 ------
 component DLI1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI1P0 ------
 component DLI1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI1P1 ------
 component DLI1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLI1P1C1 ------
 component DLI1P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 end component;


------ Component DLN0 ------
 component DLN0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN0C0 ------
 component DLN0C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN0C1 ------
 component DLN0C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN0P0 ------
 component DLN0P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN0P1 ------
 component DLN0P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN0P1C1 ------
 component DLN0P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN1 ------
 component DLN1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN1C0 ------
 component DLN1C0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN1C1 ------
 component DLN1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN1P0 ------
 component DLN1P0
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN1P1 ------
 component DLN1P1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DLN1P1C1 ------
 component DLN1P1C1
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component GND ------
 component GND
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF ------
 component INBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component INBUF_FF------
 component INBUF_FF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS15 ------
 component INBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS15D ------
 component INBUF_LVCMOS15D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS15U ------
 component INBUF_LVCMOS15U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component INBUF_LVCMOS12 ------
 component INBUF_LVCMOS12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS12D ------
 component INBUF_LVCMOS12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS12U ------
 component INBUF_LVCMOS12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS18 ------
 component INBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS18D ------
 component INBUF_LVCMOS18D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS18U ------
 component INBUF_LVCMOS18U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS25 ------
 component INBUF_LVCMOS25
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS25D ------
 component INBUF_LVCMOS25D
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS25U ------
 component INBUF_LVCMOS25U
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS33 ------
 component INBUF_LVCMOS33
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS33D ------
 component INBUF_LVCMOS33D
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS33U ------
 component INBUF_LVCMOS33U
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS5 ------
 component INBUF_LVCMOS5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS5D ------
 component INBUF_LVCMOS5D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_LVCMOS5U ------
 component INBUF_LVCMOS5U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


 ------ Component INBUF_LVDS ------
 component INBUF_LVDS
    generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

 end component;


------ Component INBUF_LVPECL ------
 component INBUF_LVPECL
     generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
                tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                             :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                             :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);

 end component;

------ Component INBUF_PCI ------
 component INBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INBUF_PCIX ------
 component INBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INV ------
 component INV
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MAJ3 ------
 component MAJ3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MAJ3X ------
 component MAJ3X
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MAJ3XI ------
 component MAJ3XI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MIN3 ------
 component MIN3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MIN3X ------
 component MIN3X
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MIN3XI ------
 component MIN3XI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2 ------
 component MX2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2A ------
 component MX2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2B ------
 component MX2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MX2C ------
 component MX2C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2 ------
 component NAND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2A ------
 component NAND2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2B ------
 component NAND2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3 ------
 component NAND3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3A ------
 component NAND3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3B ------
 component NAND3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3C ------
 component NAND3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2 ------
 component NOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2A ------
 component NOR2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2B ------
 component NOR2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3 ------
 component NOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3A ------
 component NOR3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3B ------
 component NOR3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3C ------
 component NOR3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1 ------
 component OA1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1A ------
 component OA1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1B ------
 component OA1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA1C ------
 component OA1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI1 ------
 component OAI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2 ------
 component OR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2A ------
 component OR2A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2B ------
 component OR2B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3 ------
 component OR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3A ------
 component OR3A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3B ------
 component OR3B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3C ------
 component OR3C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF ------
 component OUTBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_12 ------
 component OUTBUF_F_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_16 ------
 component OUTBUF_F_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_8 ------
 component OUTBUF_F_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_24 ------
 component OUTBUF_F_24
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS15 ------
 component OUTBUF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

------ Component OUTBUF_LVCMOS12 ------
 component OUTBUF_LVCMOS12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS18 ------
 component OUTBUF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS25 ------
 component OUTBUF_LVCMOS25
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS33 ------
 component OUTBUF_LVCMOS33
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component OUTBUF_LVCMOS5 ------
 component OUTBUF_LVCMOS5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


 
 ------ Component OUTBUF_LVDS ------
 component OUTBUF_LVDS
     generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

      tpd_D_PADP                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                                 :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :  in    STD_ULOGIC;
      PADP                           :  out   STD_ULOGIC;
      PADN                           :  out   STD_ULOGIC);
 end component;


------ Component OUTBUF_LVPECL ------
 component OUTBUF_LVPECL
     generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

      tpd_D_PADP                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :  in    STD_ULOGIC;
      PADP                           :  out   STD_ULOGIC;
      PADN                           :  out   STD_ULOGIC);

end component;

------ Component OUTBUF_PCI ------
 component OUTBUF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_PCIX ------
 component OUTBUF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_12 ------
 component OUTBUF_S_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_16 ------
 component OUTBUF_S_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_8 ------
 component OUTBUF_S_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_24 ------
 component OUTBUF_S_24
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF ------
 component TRIBUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_12 ------
 component TRIBUFF_F_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_12D ------
 component TRIBUFF_F_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_12U ------
 component TRIBUFF_F_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_16 ------
 component TRIBUFF_F_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_16D ------
 component TRIBUFF_F_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_16U ------
 component TRIBUFF_F_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_8 ------
 component TRIBUFF_F_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_8D ------
 component TRIBUFF_F_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_8U ------
 component TRIBUFF_F_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_24 ------
 component TRIBUFF_F_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_24D ------
 component TRIBUFF_F_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_24U ------
 component TRIBUFF_F_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS15 ------
 component TRIBUFF_LVCMOS15
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS15D ------
 component TRIBUFF_LVCMOS15D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS15U ------
 component TRIBUFF_LVCMOS15U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS12 ------
 component TRIBUFF_LVCMOS12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS12D ------
 component TRIBUFF_LVCMOS12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS12U ------
 component TRIBUFF_LVCMOS12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

------ Component TRIBUFF_LVCMOS18 ------
 component TRIBUFF_LVCMOS18
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS18D ------
 component TRIBUFF_LVCMOS18D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS18U ------
 component TRIBUFF_LVCMOS18U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS25 ------
 component TRIBUFF_LVCMOS25
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS25D ------
 component TRIBUFF_LVCMOS25D
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS25U ------
 component TRIBUFF_LVCMOS25U
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS33 ------
 component TRIBUFF_LVCMOS33
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS33D ------
 component TRIBUFF_LVCMOS33D
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS33U ------
 component TRIBUFF_LVCMOS33U
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS5 ------
 component TRIBUFF_LVCMOS5
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS5D ------
 component TRIBUFF_LVCMOS5D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_LVCMOS5U ------
 component TRIBUFF_LVCMOS5U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


component TRIBUFF_LVDS
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PADP              : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADP              : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_D_PADN              : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADN              : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PADP            : out   STD_ULOGIC;
                PADN            : out   STD_ULOGIC);
end component;


------ Component TRIBUFF_PCI ------
 component TRIBUFF_PCI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_PCIX ------
 component TRIBUFF_PCIX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_12 ------
 component TRIBUFF_S_12
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_12D ------
 component TRIBUFF_S_12D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_12U ------
 component TRIBUFF_S_12U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_16 ------
 component TRIBUFF_S_16
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_16D ------
 component TRIBUFF_S_16D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_16U ------
 component TRIBUFF_S_16U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_8 ------
 component TRIBUFF_S_8
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_8D ------
 component TRIBUFF_S_8D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_8U ------
 component TRIBUFF_S_8U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_24 ------
 component TRIBUFF_S_24
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_24D ------
 component TRIBUFF_S_24D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_24U ------
 component TRIBUFF_S_24U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

------ Component VCC ------
 component VCC
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 end component;


------ Component UJTAG ------
 component UJTAG
   generic(
      TimingChecksOn : Boolean := True;
      InstancePath   : STRING  := "*";
      Xon            : Boolean := False;
      MsgOn          : Boolean := True;

      tipd_UTDO      : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TMS       : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TDI       : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TCK       : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TRSTB     : VitalDelayType01 := (  0.0 ns,0.0 ns );

      tpd_TCK_UIREG0   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG1   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG2   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG3   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG4   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG5   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG6   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG7   : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TCK_URSTB    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRSH    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRCAP   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRUPD   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRCK    : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TCK_TDO      : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TRSTB_UIREG0 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG1 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG2 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG3 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG4 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG5 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG6 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG7 : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TRSTB_URSTB  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UDRSH  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UDRCAP : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UDRUPD : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TRSTB_TDO    : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TDI_UTDI     : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_TDI_TCK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_TDI_TCK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_TMS_TCK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_TMS_TCK_negedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_UTDO_TCK_posedge_negedge : VitalDelayType := 0.000 ns;
      tsetup_UTDO_TCK_negedge_negedge : VitalDelayType := 0.000 ns;

      thold_TDI_TCK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_TDI_TCK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_TMS_TCK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_TMS_TCK_negedge_posedge   : VitalDelayType := 0.000 ns;

      thold_UTDO_TCK_posedge_negedge  : VitalDelayType := 0.000 ns;
      thold_UTDO_TCK_negedge_negedge  : VitalDelayType := 0.000 ns;

      trecovery_TRSTB_TCK_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_TRSTB_TCK_posedge_posedge     : VitalDelayType := 0.000 ns;

      tpw_TCK_posedge   : VitalDelayType := 0.000 ns;
      tpw_TCK_negedge   : VitalDelayType := 0.000 ns;
      tpw_TRSTB_negedge : VitalDelayType := 0.000 ns);

   port(
      UTDO           :  in    STD_ULOGIC;
      TMS            :  in    STD_ULOGIC;
      TDI            :  in    STD_ULOGIC;
      TCK            :  in    STD_ULOGIC;
      TRSTB          :  in    STD_ULOGIC;
      UIREG0         :  out   STD_ULOGIC;
      UIREG1         :  out   STD_ULOGIC;
      UIREG2         :  out   STD_ULOGIC;
      UIREG3         :  out   STD_ULOGIC;
      UIREG4         :  out   STD_ULOGIC;
      UIREG5         :  out   STD_ULOGIC;
      UIREG6         :  out   STD_ULOGIC;
      UIREG7         :  out   STD_ULOGIC;
      UTDI           :  out   STD_ULOGIC;
      URSTB          :  out   STD_ULOGIC;
      UDRCK          :  out   STD_ULOGIC;
      UDRCAP         :  out   STD_ULOGIC;
      UDRSH          :  out   STD_ULOGIC;
      UDRUPD         :  out   STD_ULOGIC;
      TDO            :  out   STD_ULOGIC);

 end component;

------ Component XA1 ------
 component XA1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1A ------
 component XA1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1B ------
 component XA1B
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XA1C ------
 component XA1C
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XAI1 ------
 component XAI1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XAI1A ------
 component XAI1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR2 ------
 component XNOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR3 ------
 component XNOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XO1 ------
 component XO1
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XO1A ------
 component XO1A
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR2 ------
 component XOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR3 ------
 component XOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component ZOR3 ------
 component ZOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component ZOR3I ------
 component ZOR3I
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BUFF ------
 component BUFF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKINT ------
 component CLKINT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOIN_IB ------
 component IOIN_IB
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_YIN_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_YIN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		YIN		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOIN_IRC ------
 component IOIN_IRC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 end component;


------ Component IOIN_IRP ------
 component IOIN_IRP
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 end component;


------ Component IOIN_IREC ------
 component IOIN_IREC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_ICE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		ICE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 end component;


------ Component IOIN_IREP ------
 component IOIN_IREP
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		ICE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OB_EB ------
 component IOTRI_OB_EB
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_DOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		DOUT		: out    STD_ULOGIC;
		EOUT		: out    STD_ULOGIC);
 end component;


------ Component IOTRI_OB_ERC ------
 component IOTRI_OB_ERC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OB_ERP ------
 component IOTRI_OB_ERP
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OB_EREC ------
 component IOTRI_OB_EREC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OB_EREP ------
 component IOTRI_OB_EREP
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_ORC_EB ------
 component IOTRI_ORC_EB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_ORP_EB ------
 component IOTRI_ORP_EB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OREC_EB ------
 component IOTRI_OREC_EB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OREP_EB ------
 component IOTRI_OREP_EB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_ORC_ERC ------
 component IOTRI_ORC_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOTRI_OREC_EREC ------
 component IOTRI_OREC_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOTRI_ORP_ERP ------
 component IOTRI_ORP_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOTRI_OREP_EREP ------
 component IOTRI_OREP_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_EB ------
 component IOBI_IB_OB_EB
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_DOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		YIN		: in    STD_ULOGIC;
		DOUT		: out    STD_ULOGIC;
		EOUT		: out    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_ERC ------
 component IOBI_IB_OB_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_EREC ------
 component IOBI_IB_OB_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_ERP ------
 component IOBI_IB_OB_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_EREP ------
 component IOBI_IB_OB_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;

------ Component IOBI_IB_OD_EB ------
 component IOBI_IB_OD_EB
   generic (
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;

      tipd_DR          : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DF          : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E           : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OCLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_YIN         : VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_E_EOUT       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_YIN_Y        : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLR_DOUT     : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_OCLK_DOUT    : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_DR_OCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DR_OCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_DR_OCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DR_OCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

      tsetup_DF_OCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DF_OCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_DF_OCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DF_OCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

      trecovery_CLR_OCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_CLR_OCLK_negedge_posedge     : VitalDelayType := 0.000 ns;

      tpw_OCLK_posedge                   :  VitalDelayType := 0.000 ns;
      tpw_OCLK_negedge                   :  VitalDelayType := 0.000 ns;
      tperiod_OCLK_posedge               :  VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                    :  VitalDelayType := 0.000 ns
     );


   port (
      DR            :  in    std_ulogic;
      DF            :  in    std_ulogic;
      CLR           :  in    std_ulogic;
      E             :  in    std_ulogic;
      OCLK          :  in    std_ulogic;
      YIN           :  in    std_ulogic;
      DOUT          :  out   std_ulogic;
      EOUT          :  out   std_ulogic;
      Y             :  out   std_ulogic
     );
 end component;

------ Component IOBI_IB_ORC_EB ------
 component IOBI_IB_ORC_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OREC_EB ------
 component IOBI_IB_OREC_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_ORP_EB ------
 component IOBI_IB_ORP_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OREP_EB ------
 component IOBI_IB_OREP_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_ORC_ERC ------
 component IOBI_IB_ORC_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OREC_EREC ------
 component IOBI_IB_OREC_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_ORP_ERP ------
 component IOBI_IB_ORP_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OREP_EREP ------
 component IOBI_IB_OREP_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_OB_EB ------
 component IOBI_IRC_OB_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_OB_EB ------
 component IOBI_IREC_OB_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_OB_EB ------
 component IOBI_IRP_OB_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_OB_EB ------
 component IOBI_IREP_OB_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_OB_ERC ------
 component IOBI_IRC_OB_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_OB_ERC ------
 component IOBI_IREC_OB_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_OB_EREC ------
 component IOBI_IRC_OB_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_OB_EREC ------
 component IOBI_IREC_OB_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_OB_ERP ------
 component IOBI_IRP_OB_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_OB_ERP ------
 component IOBI_IREP_OB_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_OB_EREP ------
 component IOBI_IRP_OB_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_OB_EREP ------
 component IOBI_IREP_OB_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_ORC_EB ------
 component IOBI_IRC_ORC_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_ORC_EB ------
 component IOBI_IREC_ORC_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_OREC_EB ------
 component IOBI_IRC_OREC_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_OREC_EB ------
 component IOBI_IREC_OREC_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_ORP_EB ------
 component IOBI_IRP_ORP_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_OREP_EB ------
 component IOBI_IRP_OREP_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_ORP_EB ------
 component IOBI_IREP_ORP_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_OREP_EB ------
 component IOBI_IREP_OREP_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_ORC_ERC ------
 component IOBI_IRC_ORC_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRC_OREC_EREC ------
 component IOBI_IRC_OREC_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_ORC_ERC ------
 component IOBI_IREC_ORC_ERC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREC_OREC_EREC ------
 component IOBI_IREC_OREC_EREC
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_ORP_ERP ------
 component IOBI_IRP_ORP_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRP_OREP_EREP ------
 component IOBI_IRP_OREP_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_ORP_ERP ------
 component IOBI_IREP_ORP_ERP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IREP_OREP_EREP ------
 component IOBI_IREP_OREP_EREP
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOPAD_IN ------
 component IOPAD_IN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


component IOPADP_BI
    generic(
       TimingChecksOn : Boolean  := True;
       Xon            : Boolean  := False;
       InstancePath   : STRING   := "*";
       MsgOn          : Boolean  := True;

                tpw_D_posedge     : VitalDelayType    := 0.000 ns;
                tpw_D_negedge     : VitalDelayType    := 0.000 ns;
                tpw_E_posedge     : VitalDelayType    := 0.000 ns;
                tpw_E_negedge     : VitalDelayType    := 0.000 ns;
                tpw_PAD_negedge   : VitalDelayType    := 0.000 ns;
                tpw_PAD_posedge   : VitalDelayType    := 0.000 ns;
                tpw_N2PIN_negedge : VitalDelayType    := 0.000 ns;
                tpw_N2PIN_posedge : VitalDelayType    := 0.000 ns;

                tpd_D_PAD         : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PAD         : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_PAD_Y         : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_N2PIN_Y       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_D_Y           : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_Y           : VitalDelayType01  := (0.100 ns, 0.100 ns);

                tipd_D            : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_E            : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PAD          : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_N2PIN        : VitalDelayType01  := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                N2PIN           : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out   STD_ULOGIC);
end component;


 ------ Component IOPADP_IN ------
component IOPADP_IN
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
      tpw_N2PIN_posedge 	: VitalDelayType := 0.000 ns;
      tpw_N2PIN_negedge         : VitalDelayType := 0.000 ns;   

      tpd_PAD_Y                 :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_N2PIN_Y               :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD         	     :        VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_N2PIN       	     :        VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :        in    STD_ULOGIC;
      N2PIN                          :        in    STD_ULOGIC;
      Y                              :        out   STD_ULOGIC);

end component;


component IOPADN_BI
    generic(
       TimingChecksOn : Boolean  := True;
       Xon            : Boolean  := False;
       InstancePath   : STRING   := "*";
       MsgOn          : Boolean  := True;

                tpw_DB_posedge    : VitalDelayType    := 0.000 ns;
                tpw_DB_negedge    : VitalDelayType    := 0.000 ns;
                tpw_E_posedge     : VitalDelayType    := 0.000 ns;
                tpw_E_negedge     : VitalDelayType    := 0.000 ns;
                tpw_PAD_negedge   : VitalDelayType    := 0.000 ns;
                tpw_PAD_posedge   : VitalDelayType    := 0.000 ns;

                tpd_DB_PAD        : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PAD         : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_PAD_N2POUT    : VitalDelayType01  := (0.100 ns, 0.100 ns);

                tipd_DB           : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_E            : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PAD          : VitalDelayType01  := (0.000 ns, 0.000 ns));


    port(
                DB              : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                N2POUT          : out   STD_ULOGIC);
end component;


------ Component IOPADN_IN ------
component IOPADN_IN 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
 
      tpd_PAD_N2POUT                 :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD                       	     :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      N2POUT                         :	out   STD_ULOGIC);

end component;

------ Component IOPAD_TRI ------
 component IOPAD_TRI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge	: VitalDelayType := 0.000 ns;
		tpw_D_negedge	: VitalDelayType := 0.000 ns;
		tpw_E_posedge   : VitalDelayType := 0.000 ns;
		tpw_E_negedge	: VitalDelayType := 0.000 ns;

		tpd_D_PAD       : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

------ Component IOPADP_TRI ------
component IOPADP_TRI 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpw_E_posedge           : VitalDelayType := 0.000 ns;
      tpw_E_negedge           : VitalDelayType := 0.000 ns;
      tpw_D_posedge           : VitalDelayType := 0.000 ns;
      tpw_D_negedge           : VitalDelayType := 0.000 ns;
      
      tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);

end component;

------ Component IOPADN_TRI ------
component IOPADN_TRI 
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_DB_posedge 	    :   VitalDelayType := 0.000 ns;
      tpw_DB_negedge            :   VitalDelayType := 0.000 ns;
      tpw_E_posedge 		: VitalDelayType := 0.000 ns;
      tpw_E_negedge           : VitalDelayType := 0.000 ns;

      tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
      tpd_DB_PAD                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_DB                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      DB                             :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);

end component;

------ Component IOPAD_BI ------
 component IOPAD_BI
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;
  
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component IOPAD_IN_U ------
 component IOPAD_IN_U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_PAD_posedge		: VitalDelayType := 0.000 ns;
		tpw_PAD_negedge		: VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_IN_D ------
 component IOPAD_IN_D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_PAD_posedge		: VitalDelayType := 0.000 ns;
		tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_TRI_U ------
 component IOPAD_TRI_U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge	: VitalDelayType := 0.000 ns;
		tpw_D_negedge	: VitalDelayType := 0.000 ns;
		tpw_E_posedge	: VitalDelayType := 0.000 ns;
		tpw_E_negedge       : VitalDelayType := 0.000 ns;
		
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_TRI_D ------
 component IOPAD_TRI_D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge	: VitalDelayType := 0.000 ns;
	        tpw_D_negedge   : VitalDelayType := 0.000 ns;
		tpw_E_posedge   : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	: VitalDelayType := 0.000 ns;

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

------ Component IOPAD_BI_U ------
 component IOPAD_BI_U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

		tpw_D_posedge	    : VitalDelayType := 0.000 ns;
	        tpw_D_negedge       : VitalDelayType := 0.000 ns;
		tpw_E_posedge       : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_PAD_posedge     : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge     : VitalDelayType := 0.000 ns;

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);

		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOPAD_BI_D ------
 component IOPAD_BI_D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
	
		tpw_E_posedge       : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_D_posedge       : VitalDelayType := 0.000 ns;
                tpw_D_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_PAD_posedge     : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge     : VitalDelayType := 0.000 ns;

        	tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component IOPADN_OUT ------
 component IOPADN_OUT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
                tpw_DB_posedge 	: VitalDelayType := 0.000 ns;
                tpw_DB_negedge  : VitalDelayType := 0.000 ns;
		tpd_DB_PAD      : VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

------ Component BIBUF_F_2 ------
 component BIBUF_F_2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_2D ------
 component BIBUF_F_2D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_2U ------
 component BIBUF_F_2U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_4 ------
 component BIBUF_F_4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_4D ------
 component BIBUF_F_4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_4U ------
 component BIBUF_F_4U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_6 ------
 component BIBUF_F_6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_6D ------
 component BIBUF_F_6D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_F_6U ------
 component BIBUF_F_6U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_2 ------
 component BIBUF_S_2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_2D ------
 component BIBUF_S_2D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_2U ------
 component BIBUF_S_2U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_4 ------
 component BIBUF_S_4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_4D ------
 component BIBUF_S_4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_4U ------
 component BIBUF_S_4U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_6 ------
 component BIBUF_S_6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_6D ------
 component BIBUF_S_6D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BIBUF_S_6U ------
 component BIBUF_S_6U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_2 ------
 component OUTBUF_F_2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_4 ------
 component OUTBUF_F_4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_F_6 ------
 component OUTBUF_F_6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_2 ------
 component OUTBUF_S_2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_4 ------
 component OUTBUF_S_4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OUTBUF_S_6 ------
 component OUTBUF_S_6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_2 ------
 component TRIBUFF_F_2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_2D ------
 component TRIBUFF_F_2D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_2U ------
 component TRIBUFF_F_2U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_4 ------
 component TRIBUFF_F_4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_4D ------
 component TRIBUFF_F_4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_4U ------
 component TRIBUFF_F_4U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_6 ------
 component TRIBUFF_F_6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_6D ------
 component TRIBUFF_F_6D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_F_6U ------
 component TRIBUFF_F_6U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_2 ------
 component TRIBUFF_S_2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_2D ------
 component TRIBUFF_S_2D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_2U ------
 component TRIBUFF_S_2U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_4 ------
 component TRIBUFF_S_4
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_4D ------
 component TRIBUFF_S_4D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_4U ------
 component TRIBUFF_S_4U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_6 ------
 component TRIBUFF_S_6
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_6D ------
 component TRIBUFF_S_6D
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component TRIBUFF_S_6U ------
 component TRIBUFF_S_6U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component BUFD ------
 component BUFD
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INVD ------
 component INVD
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOIN_IR ------
 component IOIN_IR
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 end component;


------ Component IOIN_IRE ------
 component IOIN_IRE
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_ICE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		ICE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OB_ER ------
 component IOTRI_OB_ER
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OB_ERE ------
 component IOTRI_OB_ERE
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_OR_EB ------
 component IOTRI_OR_EB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_ORE_EB ------
 component IOTRI_ORE_EB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 end component;


------ Component IOTRI_ORE_ERE ------
 component IOTRI_ORE_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 end component;


------ Component IOTRI_OR_ER ------
 component IOTRI_OR_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_ER ------
 component IOBI_IB_OB_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OB_ERE ------
 component IOBI_IB_OB_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OR_EB ------
 component IOBI_IB_OR_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_Yin_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_Yin :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                Yin         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_ORE_EB ------
 component IOBI_IB_ORE_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_OR_ER ------
 component IOBI_IB_OR_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                YIN         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IB_ORE_ERE ------
 component IOBI_IB_ORE_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                YIN         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_OB_EB ------
 component IOBI_IR_OB_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_OB_EB ------
 component IOBI_IRE_OB_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_OB_ER ------
 component IOBI_IR_OB_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_OB_ER ------
 component IOBI_IRE_OB_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_OB_ERE ------
 component IOBI_IR_OB_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_OB_ERE ------
 component IOBI_IRE_OB_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_OR_EB ------
 component IOBI_IR_OR_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_OR_EB ------
 component IOBI_IRE_OR_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_ORE_EB ------
 component IOBI_IR_ORE_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_ORE_EB ------
 component IOBI_IRE_ORE_EB
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_OR_ER ------
 component IOBI_IR_OR_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IR_ORE_ERE ------
 component IOBI_IR_ORE_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_OR_ER ------
 component IOBI_IRE_OR_ER
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component IOBI_IRE_ORE_ERE ------
 component IOBI_IRE_ORE_ERE
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 end component;


------ Component CLKIO ------
 component CLKIO
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component CLKBIBUF ------
 component CLKBIBUF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;

------ Component PLLINT ------
component PLLINT 

    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tpd_A_Y         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                A               : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
end component;

------ Component UFROM ------
component UFROM 
  generic (

        TimingChecksOn: Boolean := True;
        InstancePath  : String  := "*";
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        MEMORYFILE    : String;
        DATA_X        : Integer := 1;
        ACT_PROGFILE      : String  := "";

        tipd_ADDR0    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR1    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR2    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR3    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR4    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR5    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR6    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_CLK      : VitalDelayType01 := ( 0.000 ns, 0.000 ns );

        tpd_CLK_DO7   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO6   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO5   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO4   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO3   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO2   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO1   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO0   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );

        tsetup_ADDR6_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR6_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR5_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR5_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR4_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR4_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR3_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR3_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR2_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR2_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR1_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR1_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR0_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR0_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tpw_CLK_posedge                   : VitalDelayType := 0.000 ns;
        tpw_CLK_negedge                   : VitalDelayType := 0.000 ns
       );

  port (
        DO0   :  out Std_ulogic := 'X';
        DO1   :  out Std_ulogic := 'X';
        DO2   :  out Std_ulogic := 'X';
        DO3   :  out Std_ulogic := 'X';
        DO4   :  out Std_ulogic := 'X';
        DO5   :  out Std_ulogic := 'X';
        DO6   :  out Std_ulogic := 'X';
        DO7   :  out Std_ulogic := 'X';
        ADDR0 :  in  Std_ulogic := 'X';
        ADDR1 :  in  Std_ulogic := 'X';
        ADDR2 :  in  Std_ulogic := 'X';
        ADDR3 :  in  Std_ulogic := 'X';
        ADDR4 :  in  Std_ulogic := 'X';
        ADDR5 :  in  Std_ulogic := 'X';
        ADDR6 :  in  Std_ulogic := 'X';
        CLK   :  in  Std_ulogic := 'X'
       );
end component;

------ Component UFROMH ------
component UFROMH 
  generic (

        TimingChecksOn: Boolean := True;
        InstancePath  : String  := "*";
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        MEMORYFILE    : String;
        DATA_X        : Integer := 1;
        ACT_PROGFILE      : String  := "";

        tipd_ADDR0    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR1    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR2    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR3    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR4    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR5    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR6    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_CLK      : VitalDelayType01 := ( 0.000 ns, 0.000 ns );

        tpd_CLK_DO7   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO6   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO5   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO4   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO3   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO2   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO1   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO0   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );

        tsetup_ADDR6_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR6_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR5_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR5_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR4_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR4_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR3_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR3_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR2_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR2_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR1_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR1_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR0_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR0_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tpw_CLK_posedge                   : VitalDelayType := 0.000 ns;
        tpw_CLK_negedge                   : VitalDelayType := 0.000 ns
       );

  port (
        DO0   :  out Std_ulogic := 'X';
        DO1   :  out Std_ulogic := 'X';
        DO2   :  out Std_ulogic := 'X';
        DO3   :  out Std_ulogic := 'X';
        DO4   :  out Std_ulogic := 'X';
        DO5   :  out Std_ulogic := 'X';
        DO6   :  out Std_ulogic := 'X';
        DO7   :  out Std_ulogic := 'X';
        ADDR0 :  in  Std_ulogic := 'X';
        ADDR1 :  in  Std_ulogic := 'X';
        ADDR2 :  in  Std_ulogic := 'X';
        ADDR3 :  in  Std_ulogic := 'X';
        ADDR4 :  in  Std_ulogic := 'X';
        ADDR5 :  in  Std_ulogic := 'X';
        ADDR6 :  in  Std_ulogic := 'X';
        CLK   :  in  Std_ulogic := 'X'
       );
end component;


------ Component ULSICC ------
component ULSICC 

    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tipd_LSICC          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                LSICC           : in    STD_ULOGIC);
end component;


------ Component ULSICC_INT ------
component ULSICC_INT 

    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tipd_USTDBY         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_LPENA          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                USTDBY          : in    STD_ULOGIC;
                LPENA           : in    STD_ULOGIC);
end component;

------ Component ULSICC_AUTH ------
component ULSICC_AUTH 

    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tipd_AUTHEN         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_LSICC          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                AUTHEN          : in    STD_ULOGIC;
                LSICC           : in    STD_ULOGIC);
end component;

------ Component SIMBUF ------
COMPONENT SIMBUF
    PORT(
                D         : in    STD_ULOGIC;
               PAD                : out    STD_ULOGIC);
END COMPONENT;

end COMPONENTS;

--------------------- END OF COMPONENTS PACKAGE SECTION  ----------------


library IEEE;
use IEEE.STD_LOGIC_1164.all;

use IEEE.VITAL_Timing.all;
use IEEE.VITAL_Primitives.all;

package VTABLES is

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

-- CLR_ipd, CLK_delayed, Q_zd, D, E_delayed, PRE_ipd, CLK_ipd
CONSTANT DFEG_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  x,  x,  L ),
( H,  L,  H,  H,  x,  x,  H,  x,  H ),
( H,  L,  H,  x,  H,  x,  H,  x,  H ),
( H,  L,  x,  H,  L,  x,  H,  x,  H ),
( H,  H,  x,  x,  x,  H,  x,  x,  S ),
( H,  x,  x,  x,  x,  L,  x,  x,  H ),
( H,  x,  x,  x,  x,  H,  L,  x,  S ),
( x,  L,  L,  L,  x,  H,  H,  x,  L ),
( x,  L,  L,  x,  H,  H,  H,  x,  L ),
( x,  L,  x,  L,  L,  H,  H,  x,  L ),
( U,  x,  L,  x,  x,  H,  x,  x,  L ),
( H,  x,  H,  x,  x,  U,  x,  x,  H )); 

-- CLR_ipd, CLK_delayed, T_delayed, Q_zd, CLK_ipd
CONSTANT tflipflop_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  L ),
( H,  L,  L,  H,  H,  x,  H ),
( H,  L,  H,  L,  H,  x,  H ),
( H,  H,  x,  x,  x,  x,  S ),
( H,  x,  x,  x,  L,  x,  S ),
( x,  L,  L,  L,  H,  x,  L ),
( x,  L,  H,  H,  H,  x,  L ));

-- CLR_ipd, CLK_delayed, PRE_delayed,K_delayed,J_delayed, Q_zd, CLK_ipd
CONSTANT jkflipflop_Q_tab : VitalStateTableType := (
( L,  x,  H,  x,  x,  x,  x,  x,  U ),
( L,  x,  L,  x,  x,  x,  x,  x,  L ),
( H,  L,  x,  L,  H,  x,  H,  x,  H ),
( H,  L,  x,  L,  x,  H,  H,  x,  H ),
( H,  L,  x,  x,  H,  L,  H,  x,  H ),
( H,  H,  L,  x,  x,  x,  x,  x,  S ),
( H,  x,  L,  x,  x,  x,  L,  x,  S ),
( H,  x,  H,  x,  x,  x,  x,  x,  H ),
( x,  L,  L,  H,  L,  x,  H,  x,  L ),
( x,  L,  L,  H,  x,  H,  H,  x,  L ),
( x,  L,  L,  x,  L,  L,  H,  x,  L ),
( U,  x,  L,  x,  x,  L,  x,  x,  L ),
( H,  x,  U,  x,  x,  H,  x,  x,  H ));

CONSTANT JKF2A_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  x,  L ),
( H,  L,  L,  H,  x,  H,  x,  H ),
( H,  L,  L,  x,  H,  H,  x,  H ),
( H,  L,  x,  H,  L,  H,  x,  H ),
( H,  H,  x,  x,  x,  x,  x,  S ),
( H,  x,  x,  x,  x,  L,  x,  S ),
( x,  L,  H,  L,  x,  H,  x,  L ),
( x,  L,  H,  x,  H,  H,  x,  L ),
( x,  L,  x,  L,  L,  H,  x,  L ),
( U,  x,  x,  x,  L,  x,  x,  L ));

CONSTANT JKF3A_Q_tab : VitalStateTableType := (
( L,  H,  L,  x,  H,  H,  x,  L ),
( L,  H,  x,  H,  H,  H,  x,  L ),
( L,  L,  H,  x,  x,  H,  x,  H ),
( L,  L,  x,  H,  x,  H,  x,  H ),
( L,  x,  L,  L,  H,  H,  x,  L ),
( L,  x,  H,  L,  x,  H,  x,  H ),
( H,  x,  x,  x,  H,  x,  x,  S ),
( x,  x,  x,  x,  L,  x,  x,  H ),
( x,  x,  x,  x,  H,  L,  x,  S ),
( x,  x,  x,  H,  U,  x,  x,  H ));


CONSTANT dlatch_DLE3B_Q_tab : VitalStateTableType := (
( x,  x,  x,  H,  x,  H ),   --active high preset

( H,  x,  x,  L,  x,  S ),   --latch
( x,  H,  x,  L,  x,  S ),   --latch

( L,  L,  H,  L,  x,  H ),   --transparent
( L,  L,  L,  L,  x,  L ),   --transparent

( U,  x,  H,  L,  H,  H ),   --o/p mux pessimism
( x,  U,  H,  L,  H,  H ),   --o/p mux pessimism
( U,  x,  L,  L,  L,  L ),   --o/p mux pessimism
( x,  U,  L,  L,  L,  L ),   --o/p mux pessimism

( L,  L,  H,  U,  x,  H ),   --PRE==X
( H,  x,  x,  U,  H,  H ),   --PRE==X
( x,  H,  x,  U,  H,  H ),   --PRE==X
( L,  U,  H,  U,  H,  H ),   --PRE==X
( U,  L,  H,  U,  H,  H ),   --PRE==X
( U,  U,  H,  U,  H,  H ));  --PRE==X
--G, E, D, P, Qn, Qn+1

CONSTANT dlatch_DLE2B_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  L ),   --active low clear

( H,  H,  x,  x,  x,  S ),   --latch
( H,  x,  H,  x,  x,  S ),   --latch

( H,  L,  L,  H,  x,  H ),   --transparent
( H,  L,  L,  L,  x,  L ),   --transparent

( H,  x,  x,  L,  L,  L ),   --o/p mux pessimism
( H,  x,  x,  H,  H,  H ),   --o/p mux pessimism

( U,  x,  x,  L,  L,  L ),   --CLR==X, o/p mux pessimism
( U,  H,  x,  x,  L,  L ),   --CLR==X, o/p mux pessimism, latch
( U,  x,  H,  x,  L,  L ),   --CLR==X, o/p mux pessimism, latch
( U,  L,  L,  L,  x,  L ));  --CLR==X, i/p mux pessimism
--C, G, E, D, Qn, Qn+1


CONSTANT dlatch_DL2C_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  L ),   --active low clear
( H,  x,  x,  H,  x,  H ),   --active high preset

( H,  H,  x,  L,  x,  S ),   --latch
( H,  L,  L,  L,  x,  L ),   --transparent

( U,  L,  L,  L,  x,  L ),   --CLR==U
( U,  H,  x,  L,  L,  L ),   --CLR==U
( x,  U,  L,  L,  L,  L ),   --CLR,G==U

( H,  U,  H,  x,  H,  H ),   --PRE==U/x,G==U
( H,  L,  H,  x,  x,  H ),   --PRE==U/x
( H,  H,  x,  U,  H,  H ));   --PRE==U
--CLR, G, D, PRE, Qn, Qn+1

CONSTANT DFN1C1_Q_tab : VitalStateTableType := (
-- CLR_ipd, CLK_ipd, D_ipd, State,   Q
(      '1',     '-',    '-',  '-',  '0' ),
(      '0',     '/',    '1',  '-',  '1' ),
(      '-',     '/',    '0',  '-',  '0' ),
(      '0',     '/',    'X',  '-',  'X' ),
(      '-',     '/',    '0',  '0',  '0' ),
(      'X',     '/',    'X',  '-',  'X' ),
(      'X',     '/',    '1',  '-',  'X' ),
(      'X',     '-',    '-',  '0',  '0' ),
(      '0',     '-',    '-',  '-',  'S' ));

end VTABLES;



--------------------- END OF VITABLE TABLE SECTION  ----------------

-- This package contains the timing for the 1.2 Volt PLL
package PLL_TIMING_V2 is
    constant EMULATED_SYSTEM_DELAY : Time := 5.700 ns; -- Delay Tap Additional CLK delay
    constant IN_DIV_DELAY          : Time := 0.850 ns; -- Input Divider intrinsic delay
    constant OUT_DIV_DELAY         : Time := 1.510 ns; -- Output Divider intrinsic delay
    constant MUX_DELAY             : Time := 1.700 ns; -- MUXA/MUXB/MUXC intrinsic delay
    constant IN_DELAY_BYP1         : Time := 1.523 ns; -- Input delay for CLKDIVDLY bypass mode - TIMING NOT UPDATED
    constant BYP_MUX_DELAY         : Time := 0.250 ns; -- Bypass MUX intrinsic delay, not used for Ys
    constant GL_DRVR_DELAY         : Time := 0.550 ns; -- Global Driver intrinsic delay
    constant Y_DRVR_DELAY          : Time := 0.000 ns; -- Y Driver intrinsic delay
    constant FB_MUX_DELAY          : Time := 1.420 ns; -- FBSEL MUX intrinsic delay
    constant X_MUX_DELAY           : Time := 0.160 ns; -- XDLYSEL MUX intrinsic delay
    constant FIN_LOCK_DELAY        : Time := 2.050 ns; -- FIN to LOCK propagation delay
    constant LOCK_OUT_DELAY        : Time := 0.820 ns; -- LOCK to OUT propagation delay
    constant PROG_INIT_DELAY       : Time := 2.300 ns;
    constant PROG_STEP_INCREMENT   : Time := 0.580 ns;
    constant BYP0_CLK_GL           : Time := 1.360 ns; -- Intrinsic delay for CLKDLY bypass mode
    constant CLKA_TO_REF_DELAY     : Time := 0.900 ns;
end PLL_TIMING_V2;

 ---- CELL AND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2 :  entity is TRUE;
 end AND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2_VITAL of AND2 is 
    for VITAL_ACT
    end for;
 end CFG_AND2_VITAL;



 ---- CELL AND2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2A :  entity is TRUE;
 end AND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2A_VITAL of AND2A is 
    for VITAL_ACT
    end for;
 end CFG_AND2A_VITAL;



 ---- CELL AND2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2B :  entity is TRUE;
 end AND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  AND  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2B_VITAL of AND2B is 
    for VITAL_ACT
    end for;
 end CFG_AND2B_VITAL;



 ---- CELL AND3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3 :  entity is TRUE;
 end AND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3_VITAL of AND3 is 
    for VITAL_ACT
    end for;
 end CFG_AND3_VITAL;



 ---- CELL AND3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3A :  entity is TRUE;
 end AND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3A_VITAL of AND3A is 
    for VITAL_ACT
    end for;
 end CFG_AND3A_VITAL;



 ---- CELL AND3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3B :  entity is TRUE;
 end AND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3B_VITAL of AND3B is 
    for VITAL_ACT
    end for;
 end CFG_AND3B_VITAL;



 ---- CELL AND3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3C :  entity is TRUE;
 end AND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AND3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3C_VITAL of AND3C is 
    for VITAL_ACT
    end for;
 end CFG_AND3C_VITAL;



 ---- CELL AO12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO12 :  entity is TRUE;
 end AO12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd ,( A_ipd  AND  (NOT B_ipd) ), (NOT C_ipd) ) OR (( (NOT A_ipd)  AND  B_ipd ) OR ( (NOT A_ipd)  AND  (NOT C_ipd) )));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO12_VITAL of AO12 is 
    for VITAL_ACT
    end for;
 end CFG_AO12_VITAL;



 ---- CELL AO13 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO13 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO13 :  entity is TRUE;
 end AO13;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO13 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR ( A_ipd  AND  (NOT C_ipd) )) OR ( B_ipd  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO13_VITAL of AO13 is 
    for VITAL_ACT
    end for;
 end CFG_AO13_VITAL;



 ---- CELL AO14 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO14 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO14 :  entity is TRUE;
 end AO14;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO14 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( (NOT A_ipd)  AND  (NOT B_ipd) ), B_ipd , C_ipd ) OR (( A_ipd  AND  B_ipd ) OR ( A_ipd  AND  (NOT C_ipd) )));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO14_VITAL of AO14 is 
    for VITAL_ACT
    end for;
 end CFG_AO14_VITAL;



 ---- CELL AO15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO15 :  entity is TRUE;
 end AO15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( A_ipd  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  (NOT B_ipd) ), C_ipd ) OR (( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO15_VITAL of AO15 is 
    for VITAL_ACT
    end for;
 end CFG_AO15_VITAL;



 ---- CELL AO16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO16 :  entity is TRUE;
 end AO16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  (NOT B_ipd) ), (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO16_VITAL of AO16 is 
    for VITAL_ACT
    end for;
 end CFG_AO16_VITAL;



 ---- CELL AO17 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO17 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO17 :  entity is TRUE;
 end AO17;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO17 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( (NOT A_ipd)  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  B_ipd ), C_ipd ) OR (( A_ipd  AND  B_ipd ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO17_VITAL of AO17 is 
    for VITAL_ACT
    end for;
 end CFG_AO17_VITAL;



 ---- CELL AO18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO18 :  entity is TRUE;
 end AO18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  B_ipd ) OR ( (NOT A_ipd)  AND  (NOT C_ipd) )) OR ( B_ipd  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO18_VITAL of AO18 is 
    for VITAL_ACT
    end for;
 end CFG_AO18_VITAL;



 ---- CELL AO1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1 :  entity is TRUE;
 end AO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1_VITAL of AO1 is 
    for VITAL_ACT
    end for;
 end CFG_AO1_VITAL;



 ---- CELL AO1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1A :  entity is TRUE;
 end AO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1A_VITAL of AO1A is 
    for VITAL_ACT
    end for;
 end CFG_AO1A_VITAL;



 ---- CELL AO1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1B :  entity is TRUE;
 end AO1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1B_VITAL of AO1B is 
    for VITAL_ACT
    end for;
 end CFG_AO1B_VITAL;



 ---- CELL AO1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1C :  entity is TRUE;
 end AO1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1C_VITAL of AO1C is 
    for VITAL_ACT
    end for;
 end CFG_AO1C_VITAL;



 ---- CELL AO1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1D :  entity is TRUE;
 end AO1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1D_VITAL of AO1D is 
    for VITAL_ACT
    end for;
 end CFG_AO1D_VITAL;



 ---- CELL AO1E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO1E is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO1E :  entity is TRUE;
 end AO1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AO1E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO1E_VITAL of AO1E is 
    for VITAL_ACT
    end for;
 end CFG_AO1E_VITAL;



 ---- CELL AOI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1 :  entity is TRUE;
 end AOI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AOI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1_VITAL of AOI1 is 
    for VITAL_ACT
    end for;
 end CFG_AOI1_VITAL;



 ---- CELL AOI1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1A :  entity is TRUE;
 end AOI1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AOI1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1A_VITAL of AOI1A is 
    for VITAL_ACT
    end for;
 end CFG_AOI1A_VITAL;



 ---- CELL AOI1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1B :  entity is TRUE;
 end AOI1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AOI1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1B_VITAL of AOI1B is 
    for VITAL_ACT
    end for;
 end CFG_AOI1B_VITAL;



 ---- CELL AOI1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1C :  entity is TRUE;
 end AOI1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AOI1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1C_VITAL of AOI1C is 
    for VITAL_ACT
    end for;
 end CFG_AOI1C_VITAL;



 ---- CELL AOI1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI1D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI1D :  entity is TRUE;
 end AOI1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AOI1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI1D_VITAL of AOI1D is 
    for VITAL_ACT
    end for;
 end CFG_AOI1D_VITAL;



 ---- CELL AOI5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI5 :  entity is TRUE;
 end AOI5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AOI5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2(( (NOT A_ipd)  AND  B_ipd ),( A_ipd  AND  (NOT B_ipd) ), C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI5_VITAL of AOI5 is 
    for VITAL_ACT
    end for;
 end CFG_AOI5_VITAL;



 ---- CELL AX1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1 :  entity is TRUE;
 end AX1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AX1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1_VITAL of AX1 is 
    for VITAL_ACT
    end for;
 end CFG_AX1_VITAL;



 ---- CELL AX1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1A :  entity is TRUE;
 end AX1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AX1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1A_VITAL of AX1A is 
    for VITAL_ACT
    end for;
 end CFG_AX1A_VITAL;



 ---- CELL AX1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1B :  entity is TRUE;
 end AX1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AX1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1B_VITAL of AX1B is 
    for VITAL_ACT
    end for;
 end CFG_AX1B_VITAL;



 ---- CELL AX1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1C :  entity is TRUE;
 end AX1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AX1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1C_VITAL of AX1C is 
    for VITAL_ACT
    end for;
 end CFG_AX1C_VITAL;



 ---- CELL AX1D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1D :  entity is TRUE;
 end AX1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AX1D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1D_VITAL of AX1D is 
    for VITAL_ACT
    end for;
 end CFG_AX1D_VITAL;



 ---- CELL AX1E ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AX1E is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AX1E :  entity is TRUE;
 end AX1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AX1E is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AX1E_VITAL of AX1E is 
    for VITAL_ACT
    end for;
 end CFG_AX1E_VITAL;



 ---- CELL AXO1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO1 :  entity is TRUE;
 end AXO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXO1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , A_ipd , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO1_VITAL of AXO1 is 
    for VITAL_ACT
    end for;
 end CFG_AXO1_VITAL;



 ---- CELL AXO2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO2 :  entity is TRUE;
 end AXO2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXO2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , (NOT A_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO2_VITAL of AXO2 is 
    for VITAL_ACT
    end for;
 end CFG_AXO2_VITAL;



 ---- CELL AXO3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO3 :  entity is TRUE;
 end AXO3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXO3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( A_ipd , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO3_VITAL of AXO3 is 
    for VITAL_ACT
    end for;
 end CFG_AXO3_VITAL;



 ---- CELL AXO5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO5 :  entity is TRUE;
 end AXO5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXO5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( B_ipd  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO5_VITAL of AXO5 is 
    for VITAL_ACT
    end for;
 end CFG_AXO5_VITAL;



 ---- CELL AXO6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO6 :  entity is TRUE;
 end AXO6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXO6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT B_ipd)  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , A_ipd , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO6_VITAL of AXO6 is 
    for VITAL_ACT
    end for;
 end CFG_AXO6_VITAL;



 ---- CELL AXO7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXO7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXO7 :  entity is TRUE;
 end AXO7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXO7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXO7_VITAL of AXO7 is 
    for VITAL_ACT
    end for;
 end CFG_AXO7_VITAL;



 ---- CELL AXOI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI1 :  entity is TRUE;
 end AXOI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXOI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , A_ipd , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI1_VITAL of AXOI1 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI1_VITAL;



 ---- CELL AXOI2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI2 :  entity is TRUE;
 end AXOI2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXOI2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  (NOT C_ipd) ) OR  VitalMUX2( C_ipd , (NOT A_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI2_VITAL of AXOI2 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI2_VITAL;



 ---- CELL AXOI3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI3 :  entity is TRUE;
 end AXOI3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXOI3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( A_ipd , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI3_VITAL of AXOI3 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI3_VITAL;



 ---- CELL AXOI4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI4 :  entity is TRUE;
 end AXOI4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXOI4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  C_ipd ) OR  VitalMUX2( A_ipd , (NOT C_ipd) , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI4_VITAL of AXOI4 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI4_VITAL;



 ---- CELL AXOI5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI5 :  entity is TRUE;
 end AXOI5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXOI5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( B_ipd  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI5_VITAL of AXOI5 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI5_VITAL;



 ---- CELL AXOI7 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AXOI7 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AXOI7 :  entity is TRUE;
 end AXOI7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of AXOI7 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT B_ipd)  AND  C_ipd ) OR  VitalMUX2( (NOT A_ipd) , (NOT C_ipd) , (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AXOI7_VITAL of AXOI7 is 
    for VITAL_ACT
    end for;
 end CFG_AXOI7_VITAL;



 ---- CELL BIBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF :  entity is TRUE;
 end BIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_VITAL of BIBUF is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_VITAL;



 ---- CELL BIBUF_F_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_12 :  entity is TRUE;
 end BIBUF_F_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_12_VITAL of BIBUF_F_12 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_12_VITAL;



 ---- CELL BIBUF_F_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_12D :  entity is TRUE;
 end BIBUF_F_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_12D_VITAL of BIBUF_F_12D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_12D_VITAL;



 ---- CELL BIBUF_F_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_12U :  entity is TRUE;
 end BIBUF_F_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_12U_VITAL of BIBUF_F_12U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_12U_VITAL;



 ---- CELL BIBUF_F_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_16 :  entity is TRUE;
 end BIBUF_F_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_16_VITAL of BIBUF_F_16 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_16_VITAL;



 ---- CELL BIBUF_F_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_16D :  entity is TRUE;
 end BIBUF_F_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_16D_VITAL of BIBUF_F_16D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_16D_VITAL;



 ---- CELL BIBUF_F_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_16U :  entity is TRUE;
 end BIBUF_F_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_16U_VITAL of BIBUF_F_16U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_16U_VITAL;



 ---- CELL BIBUF_F_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_8 :  entity is TRUE;
 end BIBUF_F_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_8_VITAL of BIBUF_F_8 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_8_VITAL;



 ---- CELL BIBUF_F_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_8D :  entity is TRUE;
 end BIBUF_F_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_8D_VITAL of BIBUF_F_8D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_8D_VITAL;



 ---- CELL BIBUF_F_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_8U :  entity is TRUE;
 end BIBUF_F_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_8U_VITAL of BIBUF_F_8U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_8U_VITAL;



 ---- CELL BIBUF_F_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_24 :  entity is TRUE;
 end BIBUF_F_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_24_VITAL of BIBUF_F_24 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_24_VITAL;



 ---- CELL BIBUF_F_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_24D :  entity is TRUE;
 end BIBUF_F_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_24D_VITAL of BIBUF_F_24D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_24D_VITAL;



 ---- CELL BIBUF_F_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_24U :  entity is TRUE;
 end BIBUF_F_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_24U_VITAL of BIBUF_F_24U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_24U_VITAL;



 ---- CELL BIBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS15 :  entity is TRUE;
 end BIBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS15_VITAL of BIBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS15_VITAL;



 ---- CELL BIBUF_LVCMOS15D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS15D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS15D :  entity is TRUE;
 end BIBUF_LVCMOS15D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS15D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS15D_VITAL of BIBUF_LVCMOS15D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS15D_VITAL;



 ---- CELL BIBUF_LVCMOS15U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS15U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS15U :  entity is TRUE;
 end BIBUF_LVCMOS15U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS15U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS15U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS15U_VITAL of BIBUF_LVCMOS15U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS15U_VITAL;


 ---- CELL BIBUF_LVCMOS12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS12 :  entity is TRUE;
 end BIBUF_LVCMOS12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS12_VITAL of BIBUF_LVCMOS12 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS12_VITAL;



 ---- CELL BIBUF_LVCMOS12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS12D :  entity is TRUE;
 end BIBUF_LVCMOS12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS12D_VITAL of BIBUF_LVCMOS12D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS12D_VITAL;



 ---- CELL BIBUF_LVCMOS12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS12U :  entity is TRUE;
 end BIBUF_LVCMOS12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS12U_VITAL of BIBUF_LVCMOS12U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS12U_VITAL;



 ---- CELL BIBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS18 :  entity is TRUE;
 end BIBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS18_VITAL of BIBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS18_VITAL;



 ---- CELL BIBUF_LVCMOS18D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS18D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS18D :  entity is TRUE;
 end BIBUF_LVCMOS18D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS18D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS18D_VITAL of BIBUF_LVCMOS18D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS18D_VITAL;



 ---- CELL BIBUF_LVCMOS18U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS18U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS18U :  entity is TRUE;
 end BIBUF_LVCMOS18U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS18U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS18U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS18U_VITAL of BIBUF_LVCMOS18U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS18U_VITAL;



 ---- CELL BIBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS25 :  entity is TRUE;
 end BIBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS25_VITAL of BIBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS25_VITAL;



 ---- CELL BIBUF_LVCMOS25D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS25D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS25D :  entity is TRUE;
 end BIBUF_LVCMOS25D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS25D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS25D_VITAL of BIBUF_LVCMOS25D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS25D_VITAL;



 ---- CELL BIBUF_LVCMOS25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS25U :  entity is TRUE;
 end BIBUF_LVCMOS25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS25U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS25U_VITAL of BIBUF_LVCMOS25U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS25U_VITAL;



 ---- CELL BIBUF_LVCMOS33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS33 is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns); 
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS33 :  entity is TRUE;
 end BIBUF_LVCMOS33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of BIBUF_LVCMOS33 is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);
        ALIAS Y_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

           -------------------------
           --  Functionality Section
           -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

          VitalPathDelay01Z (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event, tpd_E_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING,
          OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (D_ipd'last_event,tpd_D_Y, true),
                     1 => (E_ipd'last_event,tpd_E_Y, true),
                     2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS33_VITAL of BIBUF_LVCMOS33 is
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS33_VITAL;



 ---- CELL BIBUF_LVCMOS33D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS33D is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS33D :  entity is TRUE;
 end BIBUF_LVCMOS33D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of BIBUF_LVCMOS33D is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);
        ALIAS Y_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

           -------------------------
           --  Functionality Section
           -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

          VitalPathDelay01Z (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event, tpd_E_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING,
          OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (D_ipd'last_event,tpd_D_Y, true),
                     1 => (E_ipd'last_event,tpd_E_Y, true),
                     2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS33D_VITAL of BIBUF_LVCMOS33D is
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS33D_VITAL;



 ---- CELL BIBUF_LVCMOS33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS33U is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_D_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                        tpd_E_Y                 : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS33U :  entity is TRUE;
 end BIBUF_LVCMOS33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of BIBUF_LVCMOS33U is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);
        ALIAS Y_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS33U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

           -------------------------
           --  Functionality Section
           -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

          VitalPathDelay01Z (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event, tpd_E_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING,
          OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (D_ipd'last_event,tpd_D_Y, true),
                     1 => (E_ipd'last_event,tpd_E_Y, true),
                     2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;


end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS33U_VITAL of BIBUF_LVCMOS33U is
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS33U_VITAL;



 ---- CELL BIBUF_LVCMOS5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS5 :  entity is TRUE;
 end BIBUF_LVCMOS5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS5_VITAL of BIBUF_LVCMOS5 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS5_VITAL;



 ---- CELL BIBUF_LVCMOS5D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS5D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS5D :  entity is TRUE;
 end BIBUF_LVCMOS5D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS5D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS5D_VITAL of BIBUF_LVCMOS5D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS5D_VITAL;



 ---- CELL BIBUF_LVCMOS5U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVCMOS5U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVCMOS5U :  entity is TRUE;
 end BIBUF_LVCMOS5U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_LVCMOS5U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVCMOS5U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVCMOS5U_VITAL of BIBUF_LVCMOS5U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVCMOS5U_VITAL;



 ---- CELL BIBUF_LVDS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_LVDS is
    generic(
       TimingChecksOn : Boolean  := True;
       Xon            : Boolean  := False;
       InstancePath   : STRING   := "*";
       MsgOn          : Boolean  := True;

                tpw_D_posedge    : VitalDelayType    := 0.000 ns;
                tpw_D_negedge    : VitalDelayType    := 0.000 ns;
                tpw_E_posedge    : VitalDelayType    := 0.000 ns;
                tpw_E_negedge    : VitalDelayType    := 0.000 ns;
                tpw_PADP_negedge : VitalDelayType    := 0.000 ns;
                tpw_PADP_posedge : VitalDelayType    := 0.000 ns;
                tpw_PADN_negedge : VitalDelayType    := 0.000 ns;
                tpw_PADN_posedge : VitalDelayType    := 0.000 ns;

                tpd_D_PADP       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADP       : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_D_PADN       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADN       : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_PADP_Y       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_PADN_Y       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_D_Y          : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_Y          : VitalDelayType01  := (0.100 ns, 0.100 ns);

                tipd_D           : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_E           : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PADP        : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PADN        : VitalDelayType01  := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PADP            : inout STD_ULOGIC;
                PADN            : inout STD_ULOGIC;
                Y               : out   STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_LVDS :  entity is TRUE;
 end BIBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of BIBUF_LVDS is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

        SIGNAL D_ipd     : STD_ULOGIC := 'X';
        SIGNAL E_ipd     : STD_ULOGIC := 'X';
        SIGNAL PADP_ipd  : STD_ULOGIC := 'X';
        SIGNAL PADN_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
        VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd, PADP_ipd, PADN_ipd)

        -- timing check results
        VARIABLE Pviol_D         : STD_ULOGIC := '0';
        VARIABLE PeriodData_D    : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E         : STD_ULOGIC := '0';
        VARIABLE PeriodData_E    : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PADP      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PADP : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PADN      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PADN : VitalPeriodDataType := VitalPeriodDataInit;


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
        ALIAS PADP_zd    : STD_LOGIC is Results(1);
        ALIAS PADN_zd    : STD_LOGIC is Results(2);
        ALIAS Y_zd       : STD_LOGIC is Results(3);

        -- output glitch detection variables
        VARIABLE PADP_GlitchData  : VitalGlitchDataType;
        VARIABLE PADN_GlitchData  : VitalGlitchDataType;
        VARIABLE Y_GlitchData     : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PADP,
              PeriodData     => PeriodData_PADP,
              TestSignal     => PADP_ipd,
              TestSignalName => "PADP",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADP_posedge,
              PulseWidthLow  => tpw_PADP_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_PADN,
              PeriodData     => PeriodData_PADN,
              TestSignal     => PADN_ipd,
              TestSignalName => "PADN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADN_posedge,
              PulseWidthLow  => tpw_PADN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


       -------------------------
       --  Functionality Section
       -------------------------
       PADP_zd := VitalBUFIF0 (data => D_ipd, enable =>(NOT E_ipd));
       PADN_zd := VitalBUFIF0 (data => (NOT D_ipd), enable =>(NOT E_ipd));

       if ( TO_X01 ( PADP_ipd ) = '1' and TO_X01 ( PADN_ipd ) = '0' ) then
         Y_zd   := '1';
       elsif ( TO_X01 ( PADP_ipd ) = '0' and TO_X01 ( PADN_ipd ) = '1' ) then
         Y_zd   := '0';
       else
         Y_zd   := 'X';
       end if;

       ----------------------
       --  Path Delay Section
       ----------------------

       VitalPathDelay01Z (
         OutSignal     => PADP,
         GlitchData    => PADP_GlitchData,
         OutSignalName => "PADP",
         OutTemp       => PADP_zd,
         Paths    => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PADP),true),
                     1 => (E_ipd'last_event,tpd_E_PADP, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING,
         OutputMap     => "UX01ZWLH-");

       VitalPathDelay01Z (
         OutSignal     => PADN,
         GlitchData    => PADN_GlitchData,
         OutSignalName => "PADN",
         OutTemp       => PADN_zd,
         Paths    => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PADN),true),
                     1 => (E_ipd'last_event,tpd_E_PADN, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING,
         OutputMap     => "UX01ZWLH-");

       VitalPathDelay01 (
         OutSignal     => Y,
         GlitchData    => Y_GlitchData,
         OutSignalName => "Y",
         OutTemp       => Y_zd,
         Paths    => (
                     0 => (D_ipd'last_event,tpd_D_Y, true),
                     1 => (E_ipd'last_event,tpd_E_Y, true),
                     2 => (PADP_ipd'last_event,tpd_PADP_Y, true),
                     3 => (PADN_ipd'last_event,tpd_PADN_Y, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_LVDS_VITAL of BIBUF_LVDS is
    for VITAL_ACT
    end for;
 end CFG_BIBUF_LVDS_VITAL;


 ---- CELL BIBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_PCI :  entity is TRUE;
 end BIBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_PCI_VITAL of BIBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_PCI_VITAL;



 ---- CELL BIBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_PCIX :  entity is TRUE;
 end BIBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_PCIX_VITAL of BIBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_PCIX_VITAL;



 ---- CELL BIBUF_S_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_12 :  entity is TRUE;
 end BIBUF_S_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_12_VITAL of BIBUF_S_12 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_12_VITAL;



 ---- CELL BIBUF_S_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_12D :  entity is TRUE;
 end BIBUF_S_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_12D_VITAL of BIBUF_S_12D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_12D_VITAL;



 ---- CELL BIBUF_S_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_12U :  entity is TRUE;
 end BIBUF_S_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_12U_VITAL of BIBUF_S_12U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_12U_VITAL;



 ---- CELL BIBUF_S_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_16 :  entity is TRUE;
 end BIBUF_S_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_16_VITAL of BIBUF_S_16 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_16_VITAL;



 ---- CELL BIBUF_S_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_16D :  entity is TRUE;
 end BIBUF_S_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_16D_VITAL of BIBUF_S_16D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_16D_VITAL;



 ---- CELL BIBUF_S_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_16U :  entity is TRUE;
 end BIBUF_S_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_16U_VITAL of BIBUF_S_16U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_16U_VITAL;



 ---- CELL BIBUF_S_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_8 :  entity is TRUE;
 end BIBUF_S_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_8_VITAL of BIBUF_S_8 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_8_VITAL;



 ---- CELL BIBUF_S_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_8D :  entity is TRUE;
 end BIBUF_S_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_8D_VITAL of BIBUF_S_8D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_8D_VITAL;



 ---- CELL BIBUF_S_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_8U :  entity is TRUE;
 end BIBUF_S_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_8U_VITAL of BIBUF_S_8U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_8U_VITAL;



 ---- CELL BIBUF_S_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_24 :  entity is TRUE;
 end BIBUF_S_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_24_VITAL of BIBUF_S_24 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_24_VITAL;



 ---- CELL BIBUF_S_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_24D :  entity is TRUE;
 end BIBUF_S_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_24D_VITAL of BIBUF_S_24D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_24D_VITAL;



 ---- CELL BIBUF_S_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_24U :  entity is TRUE;
 end BIBUF_S_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_24U_VITAL of BIBUF_S_24U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_24U_VITAL;



 ---- CELL CLKBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF :  entity is TRUE;
 end CLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_VITAL of CLKBUF is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_VITAL;



 ---- CELL CLKBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS15 :  entity is TRUE;
 end CLKBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS15_VITAL of CLKBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS15_VITAL;


 ---- CELL CLKBUF_LVCMOS12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS12 :  entity is TRUE;
 end CLKBUF_LVCMOS12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS12_VITAL of CLKBUF_LVCMOS12 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS12_VITAL;



 ---- CELL CLKBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS18 :  entity is TRUE;
 end CLKBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS18_VITAL of CLKBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS18_VITAL;



 ---- CELL CLKBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS25 :  entity is TRUE;
 end CLKBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS25_VITAL of CLKBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS25_VITAL;



 ---- CELL CLKBUF_LVCMOS33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS33 is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS33 :  entity is TRUE;
 end CLKBUF_LVCMOS33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of CLKBUF_LVCMOS33 is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
        Y_zd :=TO_X01(PAD_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS33_VITAL of CLKBUF_LVCMOS33 is
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS33_VITAL;



 ---- CELL CLKBUF_LVCMOS5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVCMOS5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_LVCMOS5 :  entity is TRUE;
 end CLKBUF_LVCMOS5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_LVCMOS5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_LVCMOS5_VITAL of CLKBUF_LVCMOS5 is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_LVCMOS5_VITAL;



 ---- CELL CLKBUF_LVDS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBUF_LVDS : entity is TRUE;
end CLKBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

  ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)

        -- timing check results
   VARIABLE Pviol_PADP     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADP: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PADN     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADN: VitalPeriodDataType := VitalPeriodDataInit;



   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PADP,
              PeriodData     => PeriodData_PADP,
              TestSignal     => PADP_ipd,
              TestSignalName => "PADP",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADP_posedge,
              PulseWidthLow  => tpw_PADP_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_PADN,
              PeriodData     => PeriodData_PADN,
              TestSignal     => PADN_ipd,
              TestSignalName => "PADN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADN_posedge,
              PulseWidthLow  => tpw_PADN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


        end if;


      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

     ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBUF_LVDS_VITAL of CLKBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_CLKBUF_LVDS_VITAL;


 ---- CELL CLKBUF_LVPECL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;



-- entity declaration --
 entity CLKBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBUF_LVPECL : entity is TRUE;
end CLKBUF_LVPECL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)

        -- timing check results
   VARIABLE Pviol_PADP     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADP: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PADN     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADN: VitalPeriodDataType := VitalPeriodDataInit;



   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PADP,
              PeriodData     => PeriodData_PADP,
              TestSignal     => PADP_ipd,
              TestSignalName => "PADP",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADP_posedge,
              PulseWidthLow  => tpw_PADP_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVPECL",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_PADN,
              PeriodData     => PeriodData_PADN,
              TestSignal     => PADN_ipd,
              TestSignalName => "PADN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADN_posedge,
              PulseWidthLow  => tpw_PADN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_LVPECL",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


        end if;


      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBUF_LVPECL_VITAL of CLKBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_CLKBUF_LVPECL_VITAL;



 ---- CELL CLKBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_PCI :  entity is TRUE;
 end CLKBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_PCI_VITAL of CLKBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_PCI_VITAL;



 ---- CELL CLKBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBUF_PCIX :  entity is TRUE;
 end CLKBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBUF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBUF_PCIX_VITAL of CLKBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_CLKBUF_PCIX_VITAL;



 ---- CELL DFI0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0 :  entity is TRUE;
 end DFI0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFI0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed, '0', '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0_VITAL of DFI0 is
   for VITAL_ACT
   end for;
end CFG_DFI0_VITAL;



 ---- CELL DFI0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0C0 :  entity is TRUE;
 end DFI0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, QN_temp, D_delayed, '0', '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0C0_VITAL of DFI0C0 is
   for VITAL_ACT
   end for;
end CFG_DFI0C0_VITAL;



 ---- CELL DFI0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0C1 :  entity is TRUE;
 end DFI0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, QN_temp, D_delayed, '0', '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0C1_VITAL of DFI0C1 is
   for VITAL_ACT
   end for;
end CFG_DFI0C1_VITAL;



 ---- CELL DFI0E0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E0 :  entity is TRUE;
 end DFI0E0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFI0E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed, E_delayed, '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E0_VITAL of DFI0E0 is
   for VITAL_ACT
   end for;
end CFG_DFI0E0_VITAL;



 ---- CELL DFI0E0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E0C0 :  entity is TRUE;
 end DFI0E0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, QN_temp, D_delayed, E_delayed, '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E0C0_VITAL of DFI0E0C0 is
   for VITAL_ACT
   end for;
end CFG_DFI0E0C0_VITAL;



 ---- CELL DFI0E0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E0C1 :  entity is TRUE;
 end DFI0E0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, QN_temp, D_delayed, E_delayed, '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E0C1_VITAL of DFI0E0C1 is
   for VITAL_ACT
   end for;
end CFG_DFI0E0C1_VITAL;



 ---- CELL DFI0E0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E0P0 :  entity is TRUE;
 end DFI0E0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E0P0_VITAL of DFI0E0P0 is
   for VITAL_ACT
   end for;
end CFG_DFI0E0P0_VITAL;



 ---- CELL DFI0E0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E0P1 :  entity is TRUE;
 end DFI0E0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed, E_delayed, (NOT PRE_ipd), CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E0P1_VITAL of DFI0E0P1 is
   for VITAL_ACT
   end for;
end CFG_DFI0E0P1_VITAL;



 ---- CELL DFI0E1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E1 :  entity is TRUE;
 end DFI0E1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFI0E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed,  (NOT E_delayed), '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E1_VITAL of DFI0E1 is
   for VITAL_ACT
   end for;
end CFG_DFI0E1_VITAL;



 ---- CELL DFI0E1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E1C0 :  entity is TRUE;
 end DFI0E1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, QN_temp, D_delayed,  (NOT E_delayed), '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E1C0_VITAL of DFI0E1C0 is
   for VITAL_ACT
   end for;
end CFG_DFI0E1C0_VITAL;



 ---- CELL DFI0E1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E1C1 :  entity is TRUE;
 end DFI0E1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, QN_temp, D_delayed,  (NOT E_delayed), '1', CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E1C1_VITAL of DFI0E1C1 is
   for VITAL_ACT
   end for;
end CFG_DFI0E1C1_VITAL;



 ---- CELL DFI0E1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E1P0 :  entity is TRUE;
 end DFI0E1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed,  (NOT E_delayed), PRE_ipd, CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E1P0_VITAL of DFI0E1P0 is
   for VITAL_ACT
   end for;
end CFG_DFI0E1P0_VITAL;



 ---- CELL DFI0E1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0E1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0E1P1 :  entity is TRUE;
 end DFI0E1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0E1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed,  (NOT E_delayed), (NOT PRE_ipd), CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0E1P1_VITAL of DFI0E1P1 is
   for VITAL_ACT
   end for;
end CFG_DFI0E1P1_VITAL;



 ---- CELL DFI0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0P0 :  entity is TRUE;
 end DFI0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed, '0', PRE_ipd, CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0P0_VITAL of DFI0P0 is
   for VITAL_ACT
   end for;
end CFG_DFI0P0_VITAL;



 ---- CELL DFI0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0P1 :  entity is TRUE;
 end DFI0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QN_temp, D_delayed, '0', (NOT PRE_ipd), CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0P1_VITAL of DFI0P1 is
   for VITAL_ACT
   end for;
end CFG_DFI0P1_VITAL;



 ---- CELL DFI0P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI0P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI0P1C1 :  entity is TRUE;
 end DFI0P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI0P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, QN_temp, D_delayed, '0', (NOT PRE_ipd), CLK_delayed));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI0P1C1_VITAL of DFI0P1C1 is
   for VITAL_ACT
   end for;
end CFG_DFI0P1C1_VITAL;



 ---- CELL DFI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1 :  entity is TRUE;
 end DFI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFI1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed, '0', '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1_VITAL of DFI1 is
   for VITAL_ACT
   end for;
end CFG_DFI1_VITAL;



 ---- CELL DFI1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1C0 :  entity is TRUE;
 end DFI1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, QN_temp, D_delayed, '0', '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1C0_VITAL of DFI1C0 is
   for VITAL_ACT
   end for;
end CFG_DFI1C0_VITAL;



 ---- CELL DFI1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1C1 :  entity is TRUE;
 end DFI1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, QN_temp, D_delayed, '0', '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1C1_VITAL of DFI1C1 is
   for VITAL_ACT
   end for;
end CFG_DFI1C1_VITAL;



 ---- CELL DFI1E0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E0 :  entity is TRUE;
 end DFI1E0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFI1E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed, E_delayed, '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E0_VITAL of DFI1E0 is
   for VITAL_ACT
   end for;
end CFG_DFI1E0_VITAL;



 ---- CELL DFI1E0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E0C0 :  entity is TRUE;
 end DFI1E0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, QN_temp, D_delayed, E_delayed, '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E0C0_VITAL of DFI1E0C0 is
   for VITAL_ACT
   end for;
end CFG_DFI1E0C0_VITAL;



 ---- CELL DFI1E0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E0C1 :  entity is TRUE;
 end DFI1E0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, QN_temp, D_delayed, E_delayed, '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E0C1_VITAL of DFI1E0C1 is
   for VITAL_ACT
   end for;
end CFG_DFI1E0C1_VITAL;



 ---- CELL DFI1E0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E0P0 :  entity is TRUE;
 end DFI1E0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E0P0_VITAL of DFI1E0P0 is
   for VITAL_ACT
   end for;
end CFG_DFI1E0P0_VITAL;



 ---- CELL DFI1E0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E0P1 :  entity is TRUE;
 end DFI1E0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed, E_delayed, (NOT PRE_ipd), CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E0P1_VITAL of DFI1E0P1 is
   for VITAL_ACT
   end for;
end CFG_DFI1E0P1_VITAL;



 ---- CELL DFI1E1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E1 :  entity is TRUE;
 end DFI1E1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFI1E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed,  (NOT E_delayed), '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E1_VITAL of DFI1E1 is
   for VITAL_ACT
   end for;
end CFG_DFI1E1_VITAL;



 ---- CELL DFI1E1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E1C0 :  entity is TRUE;
 end DFI1E1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, QN_temp, D_delayed,  (NOT E_delayed), '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E1C0_VITAL of DFI1E1C0 is
   for VITAL_ACT
   end for;
end CFG_DFI1E1C0_VITAL;



 ---- CELL DFI1E1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E1C1 :  entity is TRUE;
 end DFI1E1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, QN_temp, D_delayed,  (NOT E_delayed), '1', CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E1C1_VITAL of DFI1E1C1 is
   for VITAL_ACT
   end for;
end CFG_DFI1E1C1_VITAL;



 ---- CELL DFI1E1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E1P0 :  entity is TRUE;
 end DFI1E1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed,  (NOT E_delayed), PRE_ipd, CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E1P0_VITAL of DFI1E1P0 is
   for VITAL_ACT
   end for;
end CFG_DFI1E1P0_VITAL;



 ---- CELL DFI1E1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1E1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1E1P1 :  entity is TRUE;
 end DFI1E1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1E1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed,  (NOT E_delayed), (NOT PRE_ipd), CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1E1P1_VITAL of DFI1E1P1 is
   for VITAL_ACT
   end for;
end CFG_DFI1E1P1_VITAL;



 ---- CELL DFI1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1P0 :  entity is TRUE;
 end DFI1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed, '0', PRE_ipd, CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1P0_VITAL of DFI1P0 is
   for VITAL_ACT
   end for;
end CFG_DFI1P0_VITAL;



 ---- CELL DFI1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1P1 :  entity is TRUE;
 end DFI1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QN_temp, D_delayed, '0', (NOT PRE_ipd), CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1P1_VITAL of DFI1P1 is
   for VITAL_ACT
   end for;
end CFG_DFI1P1_VITAL;



 ---- CELL DFI1P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFI1P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFI1P1C1 :  entity is TRUE;
 end DFI1P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFI1P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QN_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QN_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, QN_temp, D_delayed, '0', (NOT PRE_ipd), CLK_ipd));
   QN_zd := Violation XOR  (NOT QN_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_QN, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFI1P1C1_VITAL of DFI1P1C1 is
   for VITAL_ACT
   end for;
end CFG_DFI1P1C1_VITAL;



 ---- CELL DFN0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0 :  entity is TRUE;
 end DFN0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFN0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0_VITAL of DFN0 is
   for VITAL_ACT
   end for;
end CFG_DFN0_VITAL;



 ---- CELL DFN0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0C0 :  entity is TRUE;
 end DFN0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0C0_VITAL of DFN0C0 is
   for VITAL_ACT
   end for;
end CFG_DFN0C0_VITAL;



 ---- CELL DFN0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0C1 :  entity is TRUE;
 end DFN0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0C1_VITAL of DFN0C1 is
   for VITAL_ACT
   end for;
end CFG_DFN0C1_VITAL;



 ---- CELL DFN0E0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E0 :  entity is TRUE;
 end DFN0E0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFN0E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E0_VITAL of DFN0E0 is
   for VITAL_ACT
   end for;
end CFG_DFN0E0_VITAL;



 ---- CELL DFN0E0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E0C0 :  entity is TRUE;
 end DFN0E0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E0C0_VITAL of DFN0E0C0 is
   for VITAL_ACT
   end for;
end CFG_DFN0E0C0_VITAL;



 ---- CELL DFN0E0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E0C1 :  entity is TRUE;
 end DFN0E0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, Q_zd, D_delayed, E_delayed, '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E0C1_VITAL of DFN0E0C1 is
   for VITAL_ACT
   end for;
end CFG_DFN0E0C1_VITAL;



 ---- CELL DFN0E0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E0P0 :  entity is TRUE;
 end DFN0E0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN0E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E0P0_VITAL of DFN0E0P0 is
   for VITAL_ACT
   end for;
end CFG_DFN0E0P0_VITAL;



 ---- CELL DFN0E0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E0P1 :  entity is TRUE;
 end DFN0E0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN0E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, E_delayed, (NOT PRE_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E0P1_VITAL of DFN0E0P1 is
   for VITAL_ACT
   end for;
end CFG_DFN0E0P1_VITAL;



 ---- CELL DFN0E1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E1 :  entity is TRUE;
 end DFN0E1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFN0E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed,  (NOT E_delayed), '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E1_VITAL of DFN0E1 is
   for VITAL_ACT
   end for;
end CFG_DFN0E1_VITAL;



 ---- CELL DFN0E1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E1C0 :  entity is TRUE;
 end DFN0E1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_negedge,
	 Removal               => thold_CLR_CLK_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_ipd, Q_zd, D_delayed,  (NOT E_delayed), '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E1C0_VITAL of DFN0E1C0 is
   for VITAL_ACT
   end for;
end CFG_DFN0E1C0_VITAL;



 ---- CELL DFN0E1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E1C1 :  entity is TRUE;
 end DFN0E1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, Q_zd, D_delayed,  (NOT E_delayed), '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E1C1_VITAL of DFN0E1C1 is
   for VITAL_ACT
   end for;
end CFG_DFN0E1C1_VITAL;



 ---- CELL DFN0E1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E1P0 :  entity is TRUE;
 end DFN0E1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN0E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed,  (NOT E_delayed), PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E1P0_VITAL of DFN0E1P0 is
   for VITAL_ACT
   end for;
end CFG_DFN0E1P0_VITAL;



 ---- CELL DFN0E1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0E1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0E1P1 :  entity is TRUE;
 end DFN0E1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0E1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_negedge,
	 TimingData		=> Tmkr_E_CLK_negedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_negedge,
	 SetupLow		=> tsetup_E_CLK_negedge_negedge,
	 HoldHigh		=> thold_E_CLK_posedge_negedge,
	 HoldLow		=> thold_E_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN0E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_E_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed,  (NOT E_delayed), (NOT PRE_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0E1P1_VITAL of DFN0E1P1 is
   for VITAL_ACT
   end for;
end CFG_DFN0E1P1_VITAL;



 ---- CELL DFN0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0P0 :  entity is TRUE;
 end DFN0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_negedge,
	 Removal		=> thold_PRE_CLK_posedge_negedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', PRE_ipd, CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0P0_VITAL of DFN0P0 is
   for VITAL_ACT
   end for;
end CFG_DFN0P0_VITAL;



 ---- CELL DFN0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0P1 :  entity is TRUE;
 end DFN0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0P1_VITAL of DFN0P1 is
   for VITAL_ACT
   end for;
end CFG_DFN0P1_VITAL;



 ---- CELL DFN0P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN0P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN0P1C1 :  entity is TRUE;
 end DFN0P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN0P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_negedge,
	 TimingData		=> Tmkr_PRE_CLK_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_negedge,
	 Removal		=> thold_PRE_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or 
	 Tviol_PRE_CLK_negedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN0P1C1_VITAL of DFN0P1C1 is
   for VITAL_ACT
   end for;
end CFG_DFN0P1C1_VITAL;



 ---- CELL DFN1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1 :  entity is TRUE;
 end DFN1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFN1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1_VITAL of DFN1 is
   for VITAL_ACT
   end for;
end CFG_DFN1_VITAL;



 ---- CELL DFN1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1C0 :  entity is TRUE;
 end DFN1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1C0_VITAL of DFN1C0 is
   for VITAL_ACT
   end for;
end CFG_DFN1C0_VITAL;



 ---- CELL DFN1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1C1 :  entity is TRUE;
 end DFN1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 2);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFN1C1_Q_tab,
   DataIn => ( CLR_ipd, CLK_ipd, D_ipd ));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1C1_VITAL of DFN1C1 is
   for VITAL_ACT
   end for;
end CFG_DFN1C1_VITAL;



 ---- CELL DFN1E0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E0 :  entity is TRUE;
 end DFN1E0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFN1E0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E0_VITAL of DFN1E0 is
   for VITAL_ACT
   end for;
end CFG_DFN1E0_VITAL;



 ---- CELL DFN1E0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E0C0 :  entity is TRUE;
 end DFN1E0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1E0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E0C0_VITAL of DFN1E0C0 is
   for VITAL_ACT
   end for;
end CFG_DFN1E0C0_VITAL;



 ---- CELL DFN1E0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E0C1 :  entity is TRUE;
 end DFN1E0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1E0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, Q_zd, D_delayed, E_delayed, '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E0C1_VITAL of DFN1E0C1 is
   for VITAL_ACT
   end for;
end CFG_DFN1E0C1_VITAL;



 ---- CELL DFN1E0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E0P0 :  entity is TRUE;
 end DFN1E0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN1E0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, E_delayed, PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E0P0_VITAL of DFN1E0P0 is
   for VITAL_ACT
   end for;
end CFG_DFN1E0P0_VITAL;



 ---- CELL DFN1E0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E0P1 :  entity is TRUE;
 end DFN1E0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (NOT E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((NOT E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN1E0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, E_delayed, (NOT PRE_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E0P1_VITAL of DFN1E0P1 is
   for VITAL_ACT
   end for;
end CFG_DFN1E0P1_VITAL;



 ---- CELL DFN1E1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E1 :  entity is TRUE;
 end DFN1E1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "DFN1E1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed,  (NOT E_delayed), '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E1_VITAL of DFN1E1 is
   for VITAL_ACT
   end for;
end CFG_DFN1E1_VITAL;



 ---- CELL DFN1E1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E1C0 :  entity is TRUE;
 end DFN1E1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_posedge_posedge,
	 Removal               => thold_CLR_CLK_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1E1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             CLR_ipd, CLK_delayed, Q_zd, D_delayed,  (NOT E_delayed), '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E1C0_VITAL of DFN1E1C0 is
   for VITAL_ACT
   end for;
end CFG_DFN1E1C0_VITAL;



 ---- CELL DFN1E1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E1C1 :  entity is TRUE;
 end DFN1E1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1E1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, Q_zd, D_delayed,  (NOT E_delayed), '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E1C1_VITAL of DFN1E1C1 is
   for VITAL_ACT
   end for;
end CFG_DFN1E1C1_VITAL;



 ---- CELL DFN1E1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E1P0 :  entity is TRUE;
 end DFN1E1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN1E1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed,  (NOT E_delayed), PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E1P0_VITAL of DFN1E1P0 is
   for VITAL_ACT
   end for;
end CFG_DFN1E1P0_VITAL;



 ---- CELL DFN1E1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1E1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		E		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1E1P1 :  entity is TRUE;
 end DFN1E1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1E1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (E_ipd,E, tipd_E);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,E_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_E_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (E_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_CLK_posedge,
	 TimingData		=> Tmkr_E_CLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_E_CLK_posedge_posedge,
	 SetupLow		=> tsetup_E_CLK_negedge_posedge,
	 HoldHigh		=> thold_E_CLK_posedge_posedge,
	 HoldLow		=> thold_E_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((E_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN1E1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_E_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed,  (NOT E_delayed), (NOT PRE_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   E_delayed := E_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1E1P1_VITAL of DFN1E1P1 is
   for VITAL_ACT
   end for;
end CFG_DFN1E1P1_VITAL;



 ---- CELL DFN1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1P0 :  entity is TRUE;
 end DFN1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_posedge_posedge,
	 Removal		=> thold_PRE_CLK_posedge_posedge,
	 ActiveLow		 => TRUE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthLow => tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', PRE_ipd, CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1P0_VITAL of DFN1P0 is
   for VITAL_ACT
   end for;
end CFG_DFN1P0_VITAL;



 ---- CELL DFN1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1P1 :  entity is TRUE;
 end DFN1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "DFN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1P1_VITAL of DFN1P1 is
   for VITAL_ACT
   end for;
end CFG_DFN1P1_VITAL;



 ---- CELL DFN1P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFN1P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		PRE		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFN1P1C1 :  entity is TRUE;
 end DFN1P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DFN1P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_CLK_posedge,
	 TimingData		=> Tmkr_PRE_CLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_CLK_negedge_posedge,
	 Removal		=> thold_PRE_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "DFN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or 
	 Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, Q_zd, D_delayed, '0', (NOT PRE_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFN1P1C1_VITAL of DFN1P1C1 is
   for VITAL_ACT
   end for;
end CFG_DFN1P1C1_VITAL;



 ---- CELL DLI0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI0 :  entity is TRUE;
 end DLI0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLI0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLI0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI0_VITAL of DLI0 is
   for VITAL_ACT
   end for;
end CFG_DLI0_VITAL;



 ---- CELL DLI0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI0C0 :  entity is TRUE;
 end DLI0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_posedge,
	 Removal                => thold_CLR_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLI0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,G_ipd,D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI0C0_VITAL of DLI0C0 is
   for VITAL_ACT
   end for;
end CFG_DLI0C0_VITAL;



 ---- CELL DLI0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI0C1 :  entity is TRUE;
 end DLI0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLI0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),G_ipd,D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI0C1_VITAL of DLI0C1 is
   for VITAL_ACT
   end for;
end CFG_DLI0C1_VITAL;



 ---- CELL DLI0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI0P0 :  entity is TRUE;
 end DLI0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_posedge,
	 Removal                => thold_PRE_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLI0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,(NOT PRE_ipd)));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI0P0_VITAL of DLI0P0 is
   for VITAL_ACT
   end for;
end CFG_DLI0P0_VITAL;



 ---- CELL DLI0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI0P1 :  entity is TRUE;
 end DLI0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLI0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,PRE_ipd));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI0P1_VITAL of DLI0P1 is
   for VITAL_ACT
   end for;
end CFG_DLI0P1_VITAL;



 ---- CELL DLI0P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI0P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI0P1C1 :  entity is TRUE;
 end DLI0P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI0P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DLI0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),G_ipd,D_ipd,PRE_ipd));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    3 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI0P1C1_VITAL of DLI0P1C1 is
   for VITAL_ACT
   end for;
end CFG_DLI0P1C1_VITAL;



 ---- CELL DLI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI1 :  entity is TRUE;
 end DLI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLI1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLI1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI1_VITAL of DLI1 is
   for VITAL_ACT
   end for;
end CFG_DLI1_VITAL;



 ---- CELL DLI1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI1C0 :  entity is TRUE;
 end DLI1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_negedge,
	 Removal                => thold_CLR_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLI1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,(NOT G_ipd),D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI1C0_VITAL of DLI1C0 is
   for VITAL_ACT
   end for;
end CFG_DLI1C0_VITAL;



 ---- CELL DLI1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI1C1 :  entity is TRUE;
 end DLI1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_negedge,
	 Removal		=> thold_CLR_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLI1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT G_ipd),D_ipd,'0'));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI1C1_VITAL of DLI1C1 is
   for VITAL_ACT
   end for;
end CFG_DLI1C1_VITAL;



 ---- CELL DLI1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI1P0 :  entity is TRUE;
 end DLI1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_negedge,
	 Removal                => thold_PRE_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLI1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,(NOT PRE_ipd)));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI1P0_VITAL of DLI1P0 is
   for VITAL_ACT
   end for;
end CFG_DLI1P0_VITAL;



 ---- CELL DLI1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI1P1 :  entity is TRUE;
 end DLI1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_negedge,
	 Removal		=> thold_PRE_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLI1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,PRE_ipd));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI1P1_VITAL of DLI1P1 is
   for VITAL_ACT
   end for;
end CFG_DLI1P1_VITAL;



 ---- CELL DLI1P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLI1P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QN		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		QN		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLI1P1C1 :  entity is TRUE;
 end DLI1P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLI1P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QN_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QN_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QN_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_negedge,
	 Removal		=> thold_CLR_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_negedge,
	 Removal		=> thold_PRE_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DLI1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => QN_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT G_ipd),D_ipd,PRE_ipd));
	 QN_zd := Violation XOR NOT QN_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QN,
	 GlitchData => QN_GlitchData,
	 OutSignalName => "QN",
	 OutTemp => QN_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QN, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_QN, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_QN, true),
		    3 => (G_ipd'last_event, tpd_G_QN, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLI1P1C1_VITAL of DLI1P1C1 is
   for VITAL_ACT
   end for;
end CFG_DLI1P1C1_VITAL;



 ---- CELL DLN0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN0 :  entity is TRUE;
 end DLN0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLN0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLN0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN0_VITAL of DLN0 is
   for VITAL_ACT
   end for;
end CFG_DLN0_VITAL;



 ---- CELL DLN0C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN0C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN0C0 :  entity is TRUE;
 end DLN0C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN0C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_posedge,
	 Removal                => thold_CLR_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLN0C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,G_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN0C0_VITAL of DLN0C0 is
   for VITAL_ACT
   end for;
end CFG_DLN0C0_VITAL;



 ---- CELL DLN0C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN0C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN0C1 :  entity is TRUE;
 end DLN0C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN0C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLN0C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),G_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN0C1_VITAL of DLN0C1 is
   for VITAL_ACT
   end for;
end CFG_DLN0C1_VITAL;



 ---- CELL DLN0P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN0P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN0P0 :  entity is TRUE;
 end DLN0P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN0P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_posedge,
	 Removal                => thold_PRE_G_posedge_posedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLN0P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,(NOT PRE_ipd)));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN0P0_VITAL of DLN0P0 is
   for VITAL_ACT
   end for;
end CFG_DLN0P0_VITAL;



 ---- CELL DLN0P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN0P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN0P1 :  entity is TRUE;
 end DLN0P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN0P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLN0P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',G_ipd,D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN0P1_VITAL of DLN0P1 is
   for VITAL_ACT
   end for;
end CFG_DLN0P1_VITAL;



 ---- CELL DLN0P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN0P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_posedge		:  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_negedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN0P1C1 :  entity is TRUE;
 end DLN0P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN0P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_posedge,
	 TimingData		=> Tmkr_D_G_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_posedge,
	 SetupLow		=> tsetup_D_G_negedge_posedge,
	 HoldHigh		=> thold_D_G_posedge_posedge,
	 HoldLow		=> thold_D_G_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DLN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_posedge,
	 TimingData		=> Tmkr_CLR_G_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_posedge,
	 Removal		=> thold_CLR_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_posedge,
	 TimingData		=> Tmkr_PRE_G_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_posedge,
	 Removal		=> thold_PRE_G_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DLN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_G_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DLN0P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or 
		       Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),G_ipd,D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN0P1C1_VITAL of DLN0P1C1 is
   for VITAL_ACT
   end for;
end CFG_DLN0P1C1_VITAL;



 ---- CELL DLN1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN1 :  entity is TRUE;
 end DLN1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLN1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TRUE, 
	 HeaderMsg		=> InstancePath & "DLN1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN1_VITAL of DLN1 is
   for VITAL_ACT
   end for;
end CFG_DLN1_VITAL;



 ---- CELL DLN1C0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN1C0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN1C0 :  entity is TRUE;
 end DLN1C0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN1C0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_posedge_negedge,
	 Removal                => thold_CLR_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_CLR_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLN1C0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		CLR_ipd,(NOT G_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN1C0_VITAL of DLN1C0 is
   for VITAL_ACT
   end for;
end CFG_DLN1C0_VITAL;



 ---- CELL DLN1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN1C1 :  entity is TRUE;
 end DLN1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_negedge,
	 Removal		=> thold_CLR_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLN1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT G_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN1C1_VITAL of DLN1C1 is
   for VITAL_ACT
   end for;
end CFG_DLN1C1_VITAL;



 ---- CELL DLN1P0 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN1P0 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_negedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN1P0 :  entity is TRUE;
 end DLN1P0;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN1P0 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_posedge_negedge,
	 Removal                => thold_PRE_G_posedge_negedge,
	 ActiveLow		=> TRUE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthLow		=> tpw_PRE_negedge,
	 PulseWidthHigh		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLN1P0",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,(NOT PRE_ipd)));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN1P0_VITAL of DLN1P0 is
   for VITAL_ACT
   end for;
end CFG_DLN1P0_VITAL;



 ---- CELL DLN1P1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN1P1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN1P1 :  entity is TRUE;
 end DLN1P1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN1P1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_negedge,
	 Removal		=> thold_PRE_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TRUE,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	TRUE,
	 HeaderMsg		=> InstancePath & "DLN1P1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT G_ipd),D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN1P1_VITAL of DLN1P1 is
   for VITAL_ACT
   end for;
end CFG_DLN1P1_VITAL;



 ---- CELL DLN1P1C1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DLN1P1C1 is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_G_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_G_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_G_negedge		:VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_G_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_G		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		PRE		:  in    STD_ULOGIC;
		G		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DLN1P1C1 :  entity is TRUE;
 end DLN1P1C1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DLN1P1C1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL G_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (G_ipd,G, tipd_G);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, PRE_ipd,CLR_ipd,G_ipd)

	-- timing check results
	VARIABLE Tviol_D_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_G_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_G_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_G_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_G	: STD_ULOGIC := '0';
	VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_G_negedge,
	 TimingData		=> Tmkr_D_G_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_G_posedge_negedge,
	 SetupLow		=> tsetup_D_G_negedge_negedge,
	 HoldHigh		=> thold_D_G_posedge_negedge,
	 HoldLow		=> thold_D_G_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (PRE_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DLN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_G_negedge,
	 TimingData		=> Tmkr_CLR_G_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_G_negedge_negedge,
	 Removal		=> thold_CLR_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT PRE_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_PRE_G_negedge,
	 TimingData		=> Tmkr_PRE_G_negedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> G_ipd,
	 RefSignalName		=> "G",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_G_negedge_negedge,
	 Removal		=> thold_PRE_G_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DLN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_G,
	 PeriodData		=> PInfo_G,
	 TestSignal		=> G_ipd,
	 TestSignalName		=> "G",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_G_negedge,
	 PulseWidthHigh		=> tpw_G_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT PRE_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "DLN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "DLN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DLN1P1C1",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or 
		       Pviol_CLR or Pviol_G;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT G_ipd),D_ipd,PRE_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (PRE_ipd'last_event, tpd_PRE_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (G_ipd'last_event, tpd_G_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DLN1P1C1_VITAL of DLN1P1C1 is
   for VITAL_ACT
   end for;
end CFG_DLN1P1C1_VITAL;



 ---- CELL GND ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GND is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GND :  entity is TRUE;
 end GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of GND is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        Y<= '0';


end VITAL_ACT;

 configuration CFG_GND_VITAL of GND is 
    for VITAL_ACT
    end for;
 end CFG_GND_VITAL;



 ---- CELL INBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF :  entity is TRUE;
 end INBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_VITAL of INBUF is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_VITAL;


 ---- CELL INBUF_FF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_FF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_FF :  entity is TRUE;
 end INBUF_FF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_FF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_FF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_FF_VITAL of INBUF_FF is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_FF_VITAL;



 ---- CELL INBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS15 :  entity is TRUE;
 end INBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS15_VITAL of INBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS15_VITAL;



 ---- CELL INBUF_LVCMOS15D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS15D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS15D :  entity is TRUE;
 end INBUF_LVCMOS15D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS15D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS15D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS15D_VITAL of INBUF_LVCMOS15D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS15D_VITAL;



 ---- CELL INBUF_LVCMOS15U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS15U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS15U :  entity is TRUE;
 end INBUF_LVCMOS15U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS15U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS15U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS15U_VITAL of INBUF_LVCMOS15U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS15U_VITAL;


 ---- CELL INBUF_LVCMOS12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS12 :  entity is TRUE;
 end INBUF_LVCMOS12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS12_VITAL of INBUF_LVCMOS12 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS12_VITAL;



 ---- CELL INBUF_LVCMOS12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS12D :  entity is TRUE;
 end INBUF_LVCMOS12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS12D_VITAL of INBUF_LVCMOS12D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS12D_VITAL;



 ---- CELL INBUF_LVCMOS12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS12U :  entity is TRUE;
 end INBUF_LVCMOS12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS12U_VITAL of INBUF_LVCMOS12U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS12U_VITAL;



 ---- CELL INBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS18 :  entity is TRUE;
 end INBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS18_VITAL of INBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS18_VITAL;



 ---- CELL INBUF_LVCMOS18D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS18D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS18D :  entity is TRUE;
 end INBUF_LVCMOS18D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS18D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS18D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS18D_VITAL of INBUF_LVCMOS18D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS18D_VITAL;



 ---- CELL INBUF_LVCMOS18U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS18U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS18U :  entity is TRUE;
 end INBUF_LVCMOS18U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS18U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS18U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS18U_VITAL of INBUF_LVCMOS18U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS18U_VITAL;



 ---- CELL INBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS25 :  entity is TRUE;
 end INBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS25_VITAL of INBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS25_VITAL;



 ---- CELL INBUF_LVCMOS25D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS25D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS25D :  entity is TRUE;
 end INBUF_LVCMOS25D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS25D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS25D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS25D_VITAL of INBUF_LVCMOS25D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS25D_VITAL;



 ---- CELL INBUF_LVCMOS25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS25U :  entity is TRUE;
 end INBUF_LVCMOS25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS25U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS25U_VITAL of INBUF_LVCMOS25U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS25U_VITAL;



 ---- CELL INBUF_LVCMOS33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS33 is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS33 :  entity is TRUE;
 end INBUF_LVCMOS33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of INBUF_LVCMOS33 is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
        Y_zd :=TO_X01(PAD_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS33_VITAL of INBUF_LVCMOS33 is
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS33_VITAL;



 ---- CELL INBUF_LVCMOS33D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS33D is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS33D :  entity is TRUE;
 end INBUF_LVCMOS33D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of INBUF_LVCMOS33D is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS33D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS33D_VITAL of INBUF_LVCMOS33D is
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS33D_VITAL;



 ---- CELL INBUF_LVCMOS33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS33U is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_PAD_Y               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_PAD                : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                PAD             : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS33U :  entity is TRUE;
 end INBUF_LVCMOS33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of INBUF_LVCMOS33U is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS33U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS33U_VITAL of INBUF_LVCMOS33U is
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS33U_VITAL;



 ---- CELL INBUF_LVCMOS5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS5 :  entity is TRUE;
 end INBUF_LVCMOS5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS5_VITAL of INBUF_LVCMOS5 is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS5_VITAL;



 ---- CELL INBUF_LVCMOS5D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS5D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS5D :  entity is TRUE;
 end INBUF_LVCMOS5D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS5D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS5D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS5D_VITAL of INBUF_LVCMOS5D is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS5D_VITAL;



 ---- CELL INBUF_LVCMOS5U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_LVCMOS5U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_LVCMOS5U :  entity is TRUE;
 end INBUF_LVCMOS5U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_LVCMOS5U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVCMOS5U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_LVCMOS5U_VITAL of INBUF_LVCMOS5U is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_LVCMOS5U_VITAL;



  ---- CELL INBUF_LVDS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;


-- entity declaration --
 entity INBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INBUF_LVDS : entity is TRUE;
end INBUF_LVDS;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of INBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)

        -- timing check results
   VARIABLE Pviol_PADP     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADP: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PADN     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADN: VitalPeriodDataType := VitalPeriodDataInit;



  -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PADP,
              PeriodData     => PeriodData_PADP,
              TestSignal     => PADP_ipd,
              TestSignalName => "PADP",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADP_posedge,
              PulseWidthLow  => tpw_PADP_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_PADN,
              PeriodData     => PeriodData_PADN,
              TestSignal     => PADN_ipd,
              TestSignalName => "PADN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADN_posedge,
              PulseWidthLow  => tpw_PADN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


        end if;


      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

     ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INBUF_LVDS_VITAL of INBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_INBUF_LVDS_VITAL;


--   CELL INBUF_LVPECL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 -- entity declaration --
 entity INBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

      tpw_PADP_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADP_negedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_posedge        : VitalDelayType := 0.000 ns;
      tpw_PADN_negedge        : VitalDelayType := 0.000 ns;

      tpd_PADP_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_PADN_Y                    :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PADP                     :  VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PADN                     :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PADP                           :  in    STD_ULOGIC;
      PADN                           :  in    STD_ULOGIC;
      Y                              :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INBUF_LVPECL : entity is TRUE;
end INBUF_LVPECL;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of INBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PADP_ipd      : STD_ULOGIC := 'X';
   SIGNAL PADN_ipd      : STD_ULOGIC := 'X';

begin
  ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PADP_ipd, PADP, tipd_PADP);
   VitalWireDelay (PADN_ipd, PADN, tipd_PADN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PADP_ipd, PADN_ipd)

        -- timing check results
   VARIABLE Pviol_PADP     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADP: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PADN     : STD_ULOGIC := '0';
   VARIABLE PeriodData_PADN: VitalPeriodDataType := VitalPeriodDataInit;



  -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData        : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PADP,
              PeriodData     => PeriodData_PADP,
              TestSignal     => PADP_ipd,
              TestSignalName => "PADP",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADP_posedge,
              PulseWidthLow  => tpw_PADP_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVPECL",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_PADN,
              PeriodData     => PeriodData_PADN,
              TestSignal     => PADN_ipd,
              TestSignalName => "PADN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PADN_posedge,
              PulseWidthLow  => tpw_PADN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_LVPECL",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


        end if;


      -------------------------
      --  Functionality Section
      -------------------------
      if ((TO_X01(PADP_ipd) = '1') AND (TO_X01(PADN_ipd) = '0')) then
        Y_zd := '1';
      elsif ((TO_X01(PADP_ipd) = '0') AND (TO_X01(PADN_ipd) = '1')) then
        Y_zd := '0';
      else
        Y_zd := 'X';
      end if;

   ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PADP_ipd'last_event, tpd_PADP_Y, TRUE),
                 1 => (PADN_ipd'last_event, tpd_PADN_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INBUF_LVPECL_VITAL of INBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_INBUF_LVPECL_VITAL;


 ---- CELL INBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_PCI :  entity is TRUE;
 end INBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_PCI_VITAL of INBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_PCI_VITAL;



 ---- CELL INBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INBUF_PCIX :  entity is TRUE;
 end INBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)

        -- timing check results
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/INBUF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INBUF_PCIX_VITAL of INBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_INBUF_PCIX_VITAL;



 ---- CELL INV ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INV is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INV :  entity is TRUE;
 end INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INV is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INV_VITAL of INV is 
    for VITAL_ACT
    end for;
 end CFG_INV_VITAL;



 ---- CELL MAJ3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MAJ3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MAJ3 :  entity is TRUE;
 end MAJ3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MAJ3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( A_ipd  AND  B_ipd ) OR ( B_ipd  AND  C_ipd )) OR ( A_ipd  AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MAJ3_VITAL of MAJ3 is 
    for VITAL_ACT
    end for;
 end CFG_MAJ3_VITAL;



 ---- CELL MAJ3X ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MAJ3X is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MAJ3X :  entity is TRUE;
 end MAJ3X;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MAJ3X is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  B_ipd ), (NOT C_ipd) ) OR (( A_ipd  AND  (NOT B_ipd) ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MAJ3X_VITAL of MAJ3X is 
    for VITAL_ACT
    end for;
 end CFG_MAJ3X_VITAL;



 ---- CELL MAJ3XI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MAJ3XI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MAJ3XI :  entity is TRUE;
 end MAJ3XI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MAJ3XI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  B_ipd ), (NOT C_ipd) ) OR (( A_ipd  AND  (NOT B_ipd) ) AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MAJ3XI_VITAL of MAJ3XI is 
    for VITAL_ACT
    end for;
 end CFG_MAJ3XI_VITAL;



 ---- CELL MIN3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MIN3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MIN3 :  entity is TRUE;
 end MIN3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MIN3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ((( (NOT A_ipd)  AND  (NOT B_ipd) ) OR ( (NOT A_ipd)  AND  (NOT C_ipd) )) OR ( (NOT B_ipd)  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MIN3_VITAL of MIN3 is 
    for VITAL_ACT
    end for;
 end CFG_MIN3_VITAL;



 ---- CELL MIN3X ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MIN3X is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MIN3X :  entity is TRUE;
 end MIN3X;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MIN3X is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2(( A_ipd  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  (NOT B_ipd) ), (NOT C_ipd) ) OR (( (NOT A_ipd)  AND  B_ipd ) AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MIN3X_VITAL of MIN3X is 
    for VITAL_ACT
    end for;
 end CFG_MIN3X_VITAL;



 ---- CELL MIN3XI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MIN3XI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MIN3XI :  entity is TRUE;
 end MIN3XI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MIN3XI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2(( A_ipd  AND  (NOT B_ipd) ),( (NOT A_ipd)  AND  (NOT B_ipd) ), (NOT C_ipd) ) OR (( (NOT A_ipd)  AND  B_ipd ) AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MIN3XI_VITAL of MIN3XI is 
    for VITAL_ACT
    end for;
 end CFG_MIN3XI_VITAL;



 ---- CELL MX2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2 :  entity is TRUE;
 end MX2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MX2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2_VITAL of MX2 is 
    for VITAL_ACT
    end for;
 end CFG_MX2_VITAL;



 ---- CELL MX2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2A :  entity is TRUE;
 end MX2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MX2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT A_ipd) , B_ipd , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2A_VITAL of MX2A is 
    for VITAL_ACT
    end for;
 end CFG_MX2A_VITAL;



 ---- CELL MX2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2B :  entity is TRUE;
 end MX2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MX2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , (NOT B_ipd) , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2B_VITAL of MX2B is 
    for VITAL_ACT
    end for;
 end CFG_MX2B_VITAL;



 ---- CELL MX2C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MX2C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MX2C :  entity is TRUE;
 end MX2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of MX2C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( (NOT A_ipd) , (NOT B_ipd) , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MX2C_VITAL of MX2C is 
    for VITAL_ACT
    end for;
 end CFG_MX2C_VITAL;



 ---- CELL NAND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2 :  entity is TRUE;
 end NAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2_VITAL of NAND2 is 
    for VITAL_ACT
    end for;
 end CFG_NAND2_VITAL;



 ---- CELL NAND2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2A :  entity is TRUE;
 end NAND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2A_VITAL of NAND2A is 
    for VITAL_ACT
    end for;
 end CFG_NAND2A_VITAL;



 ---- CELL NAND2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2B :  entity is TRUE;
 end NAND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  AND  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2B_VITAL of NAND2B is 
    for VITAL_ACT
    end for;
 end CFG_NAND2B_VITAL;



 ---- CELL NAND3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3 :  entity is TRUE;
 end NAND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3_VITAL of NAND3 is 
    for VITAL_ACT
    end for;
 end CFG_NAND3_VITAL;



 ---- CELL NAND3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3A :  entity is TRUE;
 end NAND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3A_VITAL of NAND3A is 
    for VITAL_ACT
    end for;
 end CFG_NAND3A_VITAL;



 ---- CELL NAND3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3B :  entity is TRUE;
 end NAND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3B_VITAL of NAND3B is 
    for VITAL_ACT
    end for;
 end CFG_NAND3B_VITAL;



 ---- CELL NAND3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3C :  entity is TRUE;
 end NAND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NAND3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3C_VITAL of NAND3C is 
    for VITAL_ACT
    end for;
 end CFG_NAND3C_VITAL;



 ---- CELL NOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2 :  entity is TRUE;
 end NOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  A_ipd  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2_VITAL of NOR2 is 
    for VITAL_ACT
    end for;
 end CFG_NOR2_VITAL;



 ---- CELL NOR2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2A :  entity is TRUE;
 end NOR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2A_VITAL of NOR2A is 
    for VITAL_ACT
    end for;
 end CFG_NOR2A_VITAL;



 ---- CELL NOR2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2B :  entity is TRUE;
 end NOR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  (NOT A_ipd)  OR  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2B_VITAL of NOR2B is 
    for VITAL_ACT
    end for;
 end CFG_NOR2B_VITAL;



 ---- CELL NOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3 :  entity is TRUE;
 end NOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3_VITAL of NOR3 is 
    for VITAL_ACT
    end for;
 end CFG_NOR3_VITAL;



 ---- CELL NOR3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3A :  entity is TRUE;
 end NOR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3A_VITAL of NOR3A is 
    for VITAL_ACT
    end for;
 end CFG_NOR3A_VITAL;



 ---- CELL NOR3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3B :  entity is TRUE;
 end NOR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3B_VITAL of NOR3B is 
    for VITAL_ACT
    end for;
 end CFG_NOR3B_VITAL;



 ---- CELL NOR3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3C :  entity is TRUE;
 end NOR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of NOR3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3C_VITAL of NOR3C is 
    for VITAL_ACT
    end for;
 end CFG_NOR3C_VITAL;



 ---- CELL OA1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1 :  entity is TRUE;
 end OA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OA1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1_VITAL of OA1 is 
    for VITAL_ACT
    end for;
 end CFG_OA1_VITAL;



 ---- CELL OA1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1A :  entity is TRUE;
 end OA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OA1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1A_VITAL of OA1A is 
    for VITAL_ACT
    end for;
 end CFG_OA1A_VITAL;



 ---- CELL OA1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1B :  entity is TRUE;
 end OA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OA1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (C_ipd, A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT C_ipd)  AND ( A_ipd  OR  B_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (C_ipd'last_event,tpd_C_Y, true),
	             1 => (A_ipd'last_event,tpd_A_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1B_VITAL of OA1B is 
    for VITAL_ACT
    end for;
 end CFG_OA1B_VITAL;



 ---- CELL OA1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA1C :  entity is TRUE;
 end OA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OA1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA1C_VITAL of OA1C is 
    for VITAL_ACT
    end for;
 end CFG_OA1C_VITAL;



 ---- CELL OAI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI1 :  entity is TRUE;
 end OAI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OAI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT ( ( A_ipd  OR  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI1_VITAL of OAI1 is 
    for VITAL_ACT
    end for;
 end CFG_OAI1_VITAL;



 ---- CELL OR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2 :  entity is TRUE;
 end OR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2_VITAL of OR2 is 
    for VITAL_ACT
    end for;
 end CFG_OR2_VITAL;



 ---- CELL OR2A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2A :  entity is TRUE;
 end OR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR2A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2A_VITAL of OR2A is 
    for VITAL_ACT
    end for;
 end CFG_OR2A_VITAL;



 ---- CELL OR2B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2B :  entity is TRUE;
 end OR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR2B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  OR  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2B_VITAL of OR2B is 
    for VITAL_ACT
    end for;
 end CFG_OR2B_VITAL;



 ---- CELL OR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3 :  entity is TRUE;
 end OR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3_VITAL of OR3 is 
    for VITAL_ACT
    end for;
 end CFG_OR3_VITAL;



 ---- CELL OR3A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3A :  entity is TRUE;
 end OR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR3A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3A_VITAL of OR3A is 
    for VITAL_ACT
    end for;
 end CFG_OR3A_VITAL;



 ---- CELL OR3B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3B :  entity is TRUE;
 end OR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR3B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3B_VITAL of OR3B is 
    for VITAL_ACT
    end for;
 end CFG_OR3B_VITAL;



 ---- CELL OR3C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3C :  entity is TRUE;
 end OR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OR3C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3C_VITAL of OR3C is 
    for VITAL_ACT
    end for;
 end CFG_OR3C_VITAL;



 ---- CELL OUTBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF :  entity is TRUE;
 end OUTBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_VITAL of OUTBUF is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_VITAL;



 ---- CELL OUTBUF_F_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_12 :  entity is TRUE;
 end OUTBUF_F_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_12_VITAL of OUTBUF_F_12 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_12_VITAL;



 ---- CELL OUTBUF_F_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_16 :  entity is TRUE;
 end OUTBUF_F_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_16_VITAL of OUTBUF_F_16 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_16_VITAL;



 ---- CELL OUTBUF_F_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_8 :  entity is TRUE;
 end OUTBUF_F_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_8_VITAL of OUTBUF_F_8 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_8_VITAL;



 ---- CELL OUTBUF_F_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_24 :  entity is TRUE;
 end OUTBUF_F_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_24_VITAL of OUTBUF_F_24 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_24_VITAL;



 ---- CELL OUTBUF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS15 :  entity is TRUE;
 end OUTBUF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS15_VITAL of OUTBUF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS15_VITAL;


 ---- CELL OUTBUF_LVCMOS12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS12 :  entity is TRUE;
 end OUTBUF_LVCMOS12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS12_VITAL of OUTBUF_LVCMOS12 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS12_VITAL;



 ---- CELL OUTBUF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS18 :  entity is TRUE;
 end OUTBUF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS18_VITAL of OUTBUF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS18_VITAL;



 ---- CELL OUTBUF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS25 :  entity is TRUE;
 end OUTBUF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS25_VITAL of OUTBUF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS25_VITAL;



 ---- CELL OUTBUF_LVCMOS33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS33 is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS33 :  entity is TRUE;
 end OUTBUF_LVCMOS33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of OUTBUF_LVCMOS33 is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
        PAD_zd :=TO_X01(D_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,tpd_D_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS33_VITAL of OUTBUF_LVCMOS33 is
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS33_VITAL;



 ---- CELL OUTBUF_LVCMOS5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_LVCMOS5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_LVCMOS5 :  entity is TRUE;
 end OUTBUF_LVCMOS5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_LVCMOS5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_LVCMOS5_VITAL of OUTBUF_LVCMOS5 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_LVCMOS5_VITAL;

 

 ---- CELL OUTBUF_L ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;



-- entity declaration --
 entity OUTBUF_LVDS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

      tpd_D_PADP                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :  in    STD_ULOGIC;
      PADP                           :  out   STD_ULOGIC;
      PADN                           :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OUTBUF_LVDS : entity is TRUE;
end OUTBUF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of OUTBUF_LVDS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;




   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PADP_zd : STD_LOGIC is Results(1);
   ALIAS PADN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PADP_GlitchData     : VitalGlitchDataType;
   VARIABLE PADN_GlitchData     : VitalGlitchDataType;

   begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

      -------------------------
      --  Functionality Section
      -------------------------
      PADP_zd := TO_X01(D_ipd);
      PADN_zd := NOT(TO_X01(D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PADP,
       GlitchData => PADP_GlitchData,
       OutSignalName => "PADP",
       OutTemp => PADP_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADP, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

      VitalPathDelay01 (
       OutSignal => PADN,
       GlitchData => PADN_GlitchData,
       OutSignalName => "PADN",
       OutTemp => PADN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OUTBUF_LVDS_VITAL of OUTBUF_LVDS is
   for VITAL_ACT
   end for;
end CFG_OUTBUF_LVDS_VITAL;




 ---- CELL OUTBUF_LVPECL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;



-- entity declaration --
 entity OUTBUF_LVPECL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

      tpd_D_PADP                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_D_PADN                     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :  VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :  in    STD_ULOGIC;
      PADP                           :  out   STD_ULOGIC;
      PADN                           :  out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OUTBUF_LVPECL : entity is TRUE;
end OUTBUF_LVPECL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of OUTBUF_LVPECL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;




   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PADP_zd : STD_LOGIC is Results(1);
   ALIAS PADN_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PADP_GlitchData     : VitalGlitchDataType;
   VARIABLE PADN_GlitchData     : VitalGlitchDataType;

   begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_LVPECL",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;

      -------------------------
      --  Functionality Section
      -------------------------
      PADP_zd := TO_X01(D_ipd);
      PADN_zd := NOT(TO_X01(D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PADP,
       GlitchData => PADP_GlitchData,
       OutSignalName => "PADP",
       OutTemp => PADP_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADP, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);


      VitalPathDelay01 (
       OutSignal => PADN,
       GlitchData => PADN_GlitchData,
       OutSignalName => "PADN",
       OutTemp => PADN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PADN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OUTBUF_LVPECL_VITAL of OUTBUF_LVPECL is
   for VITAL_ACT
   end for;
end CFG_OUTBUF_LVPECL_VITAL;



 ---- CELL OUTBUF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_PCI :  entity is TRUE;
 end OUTBUF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_PCI_VITAL of OUTBUF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_PCI_VITAL;



 ---- CELL OUTBUF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_PCIX :  entity is TRUE;
 end OUTBUF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_PCIX_VITAL of OUTBUF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_PCIX_VITAL;



 ---- CELL OUTBUF_S_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_12 :  entity is TRUE;
 end OUTBUF_S_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_12_VITAL of OUTBUF_S_12 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_12_VITAL;



 ---- CELL OUTBUF_S_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_16 :  entity is TRUE;
 end OUTBUF_S_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_16_VITAL of OUTBUF_S_16 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_16_VITAL;



 ---- CELL OUTBUF_S_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_8 :  entity is TRUE;
 end OUTBUF_S_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_8_VITAL of OUTBUF_S_8 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_8_VITAL;



 ---- CELL OUTBUF_S_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_24 :  entity is TRUE;
 end OUTBUF_S_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_24_VITAL of OUTBUF_S_24 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_24_VITAL;



 ---- CELL TRIBUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF :  entity is TRUE;
 end TRIBUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_VITAL of TRIBUFF is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_VITAL;



 ---- CELL TRIBUFF_F_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_12 :  entity is TRUE;
 end TRIBUFF_F_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_12_VITAL of TRIBUFF_F_12 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_12_VITAL;



 ---- CELL TRIBUFF_F_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_12D :  entity is TRUE;
 end TRIBUFF_F_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_12D_VITAL of TRIBUFF_F_12D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_12D_VITAL;



 ---- CELL TRIBUFF_F_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_12U :  entity is TRUE;
 end TRIBUFF_F_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_12U_VITAL of TRIBUFF_F_12U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_12U_VITAL;



 ---- CELL TRIBUFF_F_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_16 :  entity is TRUE;
 end TRIBUFF_F_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_16_VITAL of TRIBUFF_F_16 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_16_VITAL;



 ---- CELL TRIBUFF_F_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_16D :  entity is TRUE;
 end TRIBUFF_F_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_16D_VITAL of TRIBUFF_F_16D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_16D_VITAL;



 ---- CELL TRIBUFF_F_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_16U :  entity is TRUE;
 end TRIBUFF_F_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_16U_VITAL of TRIBUFF_F_16U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_16U_VITAL;



 ---- CELL TRIBUFF_F_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_8 :  entity is TRUE;
 end TRIBUFF_F_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_8_VITAL of TRIBUFF_F_8 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_8_VITAL;



 ---- CELL TRIBUFF_F_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_8D :  entity is TRUE;
 end TRIBUFF_F_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_8D_VITAL of TRIBUFF_F_8D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_8D_VITAL;



 ---- CELL TRIBUFF_F_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_8U :  entity is TRUE;
 end TRIBUFF_F_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_8U_VITAL of TRIBUFF_F_8U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_8U_VITAL;



 ---- CELL TRIBUFF_F_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_24 :  entity is TRUE;
 end TRIBUFF_F_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_24_VITAL of TRIBUFF_F_24 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_24_VITAL;



 ---- CELL TRIBUFF_F_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_24D :  entity is TRUE;
 end TRIBUFF_F_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_24D_VITAL of TRIBUFF_F_24D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_24D_VITAL;



 ---- CELL TRIBUFF_F_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_24U :  entity is TRUE;
 end TRIBUFF_F_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_24U_VITAL of TRIBUFF_F_24U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_24U_VITAL;



 ---- CELL TRIBUFF_LVCMOS15 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS15 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS15 :  entity is TRUE;
 end TRIBUFF_LVCMOS15;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS15 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS15",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS15_VITAL of TRIBUFF_LVCMOS15 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS15_VITAL;



 ---- CELL TRIBUFF_LVCMOS15D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS15D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS15D :  entity is TRUE;
 end TRIBUFF_LVCMOS15D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS15D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS15D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS15D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS15D_VITAL of TRIBUFF_LVCMOS15D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS15D_VITAL;



 ---- CELL TRIBUFF_LVCMOS15U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS15U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS15U :  entity is TRUE;
 end TRIBUFF_LVCMOS15U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS15U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS15U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS15U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS15U_VITAL of TRIBUFF_LVCMOS15U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS15U_VITAL;


 ---- CELL TRIBUFF_LVCMOS12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS12 :  entity is TRUE;
 end TRIBUFF_LVCMOS12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS12_VITAL of TRIBUFF_LVCMOS12 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS12_VITAL;



 ---- CELL TRIBUFF_LVCMOS12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS12D :  entity is TRUE;
 end TRIBUFF_LVCMOS12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS12D_VITAL of TRIBUFF_LVCMOS12D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS12D_VITAL;



 ---- CELL TRIBUFF_LVCMOS12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS12U :  entity is TRUE;
 end TRIBUFF_LVCMOS12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS12U_VITAL of TRIBUFF_LVCMOS12U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS12U_VITAL;



 ---- CELL TRIBUFF_LVCMOS18 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS18 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS18 :  entity is TRUE;
 end TRIBUFF_LVCMOS18;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS18 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS18",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS18_VITAL of TRIBUFF_LVCMOS18 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS18_VITAL;



 ---- CELL TRIBUFF_LVCMOS18D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS18D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS18D :  entity is TRUE;
 end TRIBUFF_LVCMOS18D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS18D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS18D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS18D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS18D_VITAL of TRIBUFF_LVCMOS18D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS18D_VITAL;



 ---- CELL TRIBUFF_LVCMOS18U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS18U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS18U :  entity is TRUE;
 end TRIBUFF_LVCMOS18U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS18U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS18U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS18U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS18U_VITAL of TRIBUFF_LVCMOS18U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS18U_VITAL;



 ---- CELL TRIBUFF_LVCMOS25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS25 :  entity is TRUE;
 end TRIBUFF_LVCMOS25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS25",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS25_VITAL of TRIBUFF_LVCMOS25 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS25_VITAL;



 ---- CELL TRIBUFF_LVCMOS25D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS25D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS25D :  entity is TRUE;
 end TRIBUFF_LVCMOS25D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS25D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS25D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS25D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS25D_VITAL of TRIBUFF_LVCMOS25D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS25D_VITAL;



 ---- CELL TRIBUFF_LVCMOS25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS25U :  entity is TRUE;
 end TRIBUFF_LVCMOS25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS25U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS25U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS25U_VITAL of TRIBUFF_LVCMOS25U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS25U_VITAL;



 ---- CELL TRIBUFF_LVCMOS33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS33 is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS33 :  entity is TRUE;
 end TRIBUFF_LVCMOS33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of TRIBUFF_LVCMOS33 is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS33",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


           ----------------------
           --  Path Delay Section
           ----------------------


          VitalPathDelay01Z (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event, tpd_E_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING,
          OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS33_VITAL of TRIBUFF_LVCMOS33 is
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS33_VITAL;



 ---- CELL TRIBUFF_LVCMOS33D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS33D is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS33D :  entity is TRUE;
 end TRIBUFF_LVCMOS33D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of TRIBUFF_LVCMOS33D is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        end block;


        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS33D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS33D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


           ----------------------
           --  Path Delay Section
           ----------------------

          VitalPathDelay01Z (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event, tpd_E_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING,
          OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS33D_VITAL of TRIBUFF_LVCMOS33D is
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS33D_VITAL;



 ---- CELL TRIBUFF_LVCMOS33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS33U is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PAD               : VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS33U :  entity is TRUE;
 end TRIBUFF_LVCMOS33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of TRIBUFF_LVCMOS33U is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS PAD_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS33U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS33U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


           -------------------------
           --  Functionality Section
           -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


           ----------------------
           --  Path Delay Section
           ----------------------

          VitalPathDelay01Z (
           OutSignal => PAD,
           GlitchData => PAD_GlitchData,
           OutSignalName => "PAD",
           OutTemp => PAD_zd,
           Paths => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event, tpd_E_PAD, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING,
          OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS33U_VITAL of TRIBUFF_LVCMOS33U is
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS33U_VITAL;



 ---- CELL TRIBUFF_LVCMOS5 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS5 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS5 :  entity is TRUE;
 end TRIBUFF_LVCMOS5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS5 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS5",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS5_VITAL of TRIBUFF_LVCMOS5 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS5_VITAL;



 ---- CELL TRIBUFF_LVCMOS5D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS5D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS5D :  entity is TRUE;
 end TRIBUFF_LVCMOS5D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS5D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS5D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS5D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS5D_VITAL of TRIBUFF_LVCMOS5D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS5D_VITAL;



 ---- CELL TRIBUFF_LVCMOS5U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVCMOS5U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVCMOS5U :  entity is TRUE;
 end TRIBUFF_LVCMOS5U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_LVCMOS5U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS5U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVCMOS5U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVCMOS5U_VITAL of TRIBUFF_LVCMOS5U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVCMOS5U_VITAL;



 ---- CELL TRIBUFF_LVDS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_LVDS is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

                tpd_D_PADP              : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADP              : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_D_PADN              : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PADN              : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tipd_D          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PADP            : out   STD_ULOGIC;
                PADN            : out   STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_LVDS :  entity is TRUE;
 end TRIBUFF_LVDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of TRIBUFF_LVDS is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (D_ipd, D, tipd_D);
        VitalWireDelay (E_ipd, E, tipd_E);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(0 to 1)  := (others => 'X');
        ALIAS PADP_zd : STD_LOGIC is Results(0);
        ALIAS PADN_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE PADP_GlitchData  : VitalGlitchDataType;
        VARIABLE PADN_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_LVDS",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


       -------------------------
       --  Functionality Section
       -------------------------

       PADP_zd := VitalBUFIF0 (data => D_ipd, enable =>(NOT E_ipd));
       PADN_zd := VitalBUFIF0 (data => (NOT D_ipd), enable =>(NOT E_ipd));

       ----------------------
       --  Path Delay Section
       ----------------------

       VitalPathDelay01Z (
         OutSignal     => PADP,
         GlitchData    => PADP_GlitchData,
         OutSignalName => "PADP",
         OutTemp       => PADP_zd,
         Paths   => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PADP),true),
                     1 => (E_ipd'last_event,tpd_E_PADP, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING,
         OutputMap     => "UX01ZWLH-");

       VitalPathDelay01Z (
         OutSignal     => PADN,
         GlitchData    => PADN_GlitchData,
         OutSignalName => "PADN",
         OutTemp       => PADN_zd,
         Paths   => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PADN),true),
                     1 => (E_ipd'last_event,tpd_E_PADN, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING,
         OutputMap     => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_LVDS_VITAL of TRIBUFF_LVDS is
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_LVDS_VITAL;



 ---- CELL TRIBUFF_PCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_PCI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_PCI :  entity is TRUE;
 end TRIBUFF_PCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_PCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_PCI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_PCI_VITAL of TRIBUFF_PCI is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_PCI_VITAL;



 ---- CELL TRIBUFF_PCIX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_PCIX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_PCIX :  entity is TRUE;
 end TRIBUFF_PCIX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_PCIX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_PCIX",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_PCIX_VITAL of TRIBUFF_PCIX is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_PCIX_VITAL;



 ---- CELL TRIBUFF_S_12 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_12 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_12 :  entity is TRUE;
 end TRIBUFF_S_12;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_12 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_12",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_12_VITAL of TRIBUFF_S_12 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_12_VITAL;



 ---- CELL TRIBUFF_S_12D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_12D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_12D :  entity is TRUE;
 end TRIBUFF_S_12D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_12D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_12D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_12D_VITAL of TRIBUFF_S_12D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_12D_VITAL;



 ---- CELL TRIBUFF_S_12U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_12U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_12U :  entity is TRUE;
 end TRIBUFF_S_12U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_12U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_12U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_12U_VITAL of TRIBUFF_S_12U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_12U_VITAL;



 ---- CELL TRIBUFF_S_16 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_16 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_16 :  entity is TRUE;
 end TRIBUFF_S_16;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_16 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_16",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_16_VITAL of TRIBUFF_S_16 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_16_VITAL;



 ---- CELL TRIBUFF_S_16D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_16D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_16D :  entity is TRUE;
 end TRIBUFF_S_16D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_16D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_16D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_16D_VITAL of TRIBUFF_S_16D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_16D_VITAL;



 ---- CELL TRIBUFF_S_16U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_16U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_16U :  entity is TRUE;
 end TRIBUFF_S_16U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_16U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_16U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_16U_VITAL of TRIBUFF_S_16U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_16U_VITAL;



 ---- CELL TRIBUFF_S_8 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_8 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_8 :  entity is TRUE;
 end TRIBUFF_S_8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_8 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_8",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_8_VITAL of TRIBUFF_S_8 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_8_VITAL;



 ---- CELL TRIBUFF_S_8D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_8D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_8D :  entity is TRUE;
 end TRIBUFF_S_8D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_8D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_8D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_8D_VITAL of TRIBUFF_S_8D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_8D_VITAL;



 ---- CELL TRIBUFF_S_8U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_8U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_8U :  entity is TRUE;
 end TRIBUFF_S_8U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_8U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_8U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_8U_VITAL of TRIBUFF_S_8U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_8U_VITAL;



 ---- CELL TRIBUFF_S_24 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_24 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_24 :  entity is TRUE;
 end TRIBUFF_S_24;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_24 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_24",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_24_VITAL of TRIBUFF_S_24 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_24_VITAL;



 ---- CELL TRIBUFF_S_24D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_24D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_24D :  entity is TRUE;
 end TRIBUFF_S_24D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_24D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_24D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_24D_VITAL of TRIBUFF_S_24D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_24D_VITAL;



 ---- CELL TRIBUFF_S_24U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_24U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_24U :  entity is TRUE;
 end TRIBUFF_S_24U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_24U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_24U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_24U_VITAL of TRIBUFF_S_24U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_24U_VITAL;



 ---- CELL VCC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity VCC is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of VCC :  entity is TRUE;
 end VCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of VCC is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        Y<= '1';


end VITAL_ACT;

 configuration CFG_VCC_VITAL of VCC is 
    for VITAL_ACT
    end for;
 end CFG_VCC_VITAL;



 ---- CELL XA1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1 :  entity is TRUE;
 end XA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XA1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1_VITAL of XA1 is 
    for VITAL_ACT
    end for;
 end CFG_XA1_VITAL;



 ---- CELL XA1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1A :  entity is TRUE;
 end XA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XA1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1A_VITAL of XA1A is 
    for VITAL_ACT
    end for;
 end CFG_XA1A_VITAL;



 ---- CELL XA1B ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1B is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1B :  entity is TRUE;
 end XA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XA1B is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1B_VITAL of XA1B is 
    for VITAL_ACT
    end for;
 end CFG_XA1B_VITAL;



 ---- CELL XA1C ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XA1C is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XA1C :  entity is TRUE;
 end XA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XA1C is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XA1C_VITAL of XA1C is 
    for VITAL_ACT
    end for;
 end CFG_XA1C_VITAL;



 ---- CELL XAI1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XAI1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XAI1 :  entity is TRUE;
 end XAI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XAI1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XAI1_VITAL of XAI1 is 
    for VITAL_ACT
    end for;
 end CFG_XAI1_VITAL;



 ---- CELL XAI1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XAI1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XAI1A :  entity is TRUE;
 end XAI1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XAI1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XAI1A_VITAL of XAI1A is 
    for VITAL_ACT
    end for;
 end CFG_XAI1A_VITAL;



 ---- CELL XNOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR2 :  entity is TRUE;
 end XNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XNOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR2_VITAL of XNOR2 is 
    for VITAL_ACT
    end for;
 end CFG_XNOR2_VITAL;



 ---- CELL XNOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR3 :  entity is TRUE;
 end XNOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XNOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT (  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR3_VITAL of XNOR3 is 
    for VITAL_ACT
    end for;
 end CFG_XNOR3_VITAL;



 ---- CELL XO1 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XO1 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XO1 :  entity is TRUE;
 end XO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XO1 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XO1_VITAL of XO1 is 
    for VITAL_ACT
    end for;
 end CFG_XO1_VITAL;



 ---- CELL XO1A ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XO1A is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XO1A :  entity is TRUE;
 end XO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XO1A is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XO1A_VITAL of XO1A is 
    for VITAL_ACT
    end for;
 end CFG_XO1A_VITAL;



 ---- CELL XOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR2 :  entity is TRUE;
 end XOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR2_VITAL of XOR2 is 
    for VITAL_ACT
    end for;
 end CFG_XOR2_VITAL;



 ---- CELL XOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR3 :  entity is TRUE;
 end XOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of XOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) ) XOR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR3_VITAL of XOR3 is 
    for VITAL_ACT
    end for;
 end CFG_XOR3_VITAL;



 ---- CELL ZOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ZOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of ZOR3 :  entity is TRUE;
 end ZOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of ZOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  (NOT B_ipd) ), C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_ZOR3_VITAL of ZOR3 is 
    for VITAL_ACT
    end for;
 end CFG_ZOR3_VITAL;



 ---- CELL ZOR3I ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity ZOR3I is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of ZOR3I :  entity is TRUE;
 end ZOR3I;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of ZOR3I is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2(( A_ipd  AND  B_ipd ),( (NOT A_ipd)  AND  (NOT B_ipd) ), C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_ZOR3I_VITAL of ZOR3I is 
    for VITAL_ACT
    end for;
 end CFG_ZOR3I_VITAL;



 ---- CELL BUFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BUFF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BUFF :  entity is TRUE;
 end BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BUFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BUFF_VITAL of BUFF is 
    for VITAL_ACT
    end for;
 end CFG_BUFF_VITAL;

 
 ---- CELL CLKINT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKINT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKINT :  entity is TRUE;
 end CLKINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKINT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKINT_VITAL of CLKINT is 
    for VITAL_ACT
    end for;
 end CFG_CLKINT_VITAL;


 ---- CELL IOIN_IB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IB is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_YIN_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_YIN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		YIN		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOIN_IB :  entity is TRUE;
 end IOIN_IB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (YIN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(YIN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (YIN_ipd'last_event,tpd_YIN_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOIN_IB_VITAL of IOIN_IB is 
    for VITAL_ACT
    end for;
 end CFG_IOIN_IB_VITAL;



 ---- CELL IOIN_IRC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IRC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_IRC :  entity is TRUE;
 end IOIN_IRC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IRC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, CLR_ipd,ICLK_ipd)

	-- timing check results
	VARIABLE Tviol_YIN_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_YIN_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_ICLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_ICLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE ICLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE YIN_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_YIN_ICLK_posedge,
	 TimingData		=> Tmkr_YIN_ICLK_posedge,
	 TestSignal		=> YIN_ipd,
	 TestSignalName		=> "YIN",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName	        => "ICLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_YIN_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_YIN_ICLK_negedge_posedge,
	 HoldHigh		=> thold_YIN_ICLK_posedge_posedge,
	 HoldLow		=> thold_YIN_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOIN_IRC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_ICLK_posedge,
	 TimingData             => Tmkr_CLR_ICLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => ICLK_ipd,
	 RefSignalName          => "ICLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_ICLK_negedge_posedge,
	 Removal               => thold_CLR_ICLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IRC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_ICLK,
	 PeriodData		=> PInfo_ICLK,
	 TestSignal		=> ICLK_ipd,
	 TestSignalName		=> "ICLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_ICLK_posedge,
	 PulseWidthLow		=> tpw_ICLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOIN_IRC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOIN_IRC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_YIN_ICLK_posedge or 
	 Pviol_CLR or 
	 Pviol_ICLK;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Y,
	 GlitchData => Y_GlitchData,
	 OutSignalName => "Y",
	 OutTemp => Y_zd,
	 Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Y, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOIN_IRC_VITAL of IOIN_IRC is
   for VITAL_ACT
   end for;
end CFG_IOIN_IRC_VITAL;



 ---- CELL IOIN_IRP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IRP is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_IRP :  entity is TRUE;
 end IOIN_IRP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IRP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, PRE_ipd,ICLK_ipd)

	-- timing check results
	VARIABLE Tviol_YIN_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_YIN_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_ICLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_ICLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE ICLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE YIN_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_YIN_ICLK_posedge,
	 TimingData		=> Tmkr_YIN_ICLK_posedge,
	 TestSignal		=> YIN_ipd,
	 TestSignalName		=> "YIN",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName	        => "ICLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_YIN_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_YIN_ICLK_negedge_posedge,
	 HoldHigh		=> thold_YIN_ICLK_posedge_posedge,
	 HoldLow		=> thold_YIN_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOIN_IRP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_ICLK_posedge,
	 TimingData		=> Tmkr_PRE_ICLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName		=> "ICLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_ICLK_negedge_posedge,
	 Removal		=> thold_PRE_ICLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IRP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_ICLK,
	 PeriodData		=> PInfo_ICLK,
	 TestSignal		=> ICLK_ipd,
	 TestSignalName		=> "ICLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_ICLK_posedge,
	 PulseWidthLow		=> tpw_ICLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOIN_IRP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "IOIN_IRP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_YIN_ICLK_posedge or 
	 Tviol_PRE_ICLK_posedge or 
	 Tviol_PRE_ICLK_posedge or Pviol_PRE or Pviol_ICLK;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Y,
	 GlitchData => Y_GlitchData,
	 OutSignalName => "Y",
	 OutTemp => Y_zd,
	 Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Y, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOIN_IRP_VITAL of IOIN_IRP is
   for VITAL_ACT
   end for;
end CFG_IOIN_IRP_VITAL;



 ---- CELL IOIN_IREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IREC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_ICE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		ICE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_IREC :  entity is TRUE;
 end IOIN_IREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IREC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (ICE_ipd,ICE, tipd_ICE);
	  VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, CLR_ipd,ICE_ipd,ICLK_ipd)

	-- timing check results
	VARIABLE Tviol_YIN_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_YIN_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_ICE_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_ICE_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_ICLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_ICLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE ICE_delayed	: STD_ULOGIC := 'X';
	VARIABLE ICLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE YIN_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_YIN_ICLK_posedge,
	 TimingData		=> Tmkr_YIN_ICLK_posedge,
	 TestSignal		=> YIN_ipd,
	 TestSignalName		=> "YIN",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName	        => "ICLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_YIN_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_YIN_ICLK_negedge_posedge,
	 HoldHigh		=> thold_YIN_ICLK_posedge_posedge,
	 HoldLow		=> thold_YIN_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (ICE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOIN_IREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_ICE_ICLK_posedge,
	 TimingData		=> Tmkr_ICE_ICLK_posedge,
	 TestSignal		=> ICE_ipd,
	 TestSignalName		=> "ICE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName		=> "ICLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_ICE_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_ICE_ICLK_negedge_posedge,
	 HoldHigh		=> thold_ICE_ICLK_posedge_posedge,
	 HoldLow		=> thold_ICE_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_ICLK_posedge,
	 TimingData             => Tmkr_CLR_ICLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => ICLK_ipd,
	 RefSignalName          => "ICLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_ICLK_negedge_posedge,
	 Removal               => thold_CLR_ICLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((ICE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_ICLK,
	 PeriodData		=> PInfo_ICLK,
	 TestSignal		=> ICLK_ipd,
	 TestSignalName		=> "ICLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_ICLK_posedge,
	 PulseWidthLow		=> tpw_ICLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOIN_IREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOIN_IREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_YIN_ICLK_posedge or 
	 Tviol_ICE_ICLK_posedge or 
	 Pviol_CLR or Pviol_ICLK;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Y,
	 GlitchData => Y_GlitchData,
	 OutSignalName => "Y",
	 OutTemp => Y_zd,
	 Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Y, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOIN_IREC_VITAL of IOIN_IREC is
   for VITAL_ACT
   end for;
end CFG_IOIN_IREC_VITAL;



 ---- CELL IOIN_IREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IREP is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		ICE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_IREP :  entity is TRUE;
 end IOIN_IREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IREP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICE_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (ICE_ipd,ICE, tipd_ICE);
	  VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, PRE_ipd,ICE_ipd,ICLK_ipd)

	-- timing check results
	VARIABLE Tviol_YIN_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_YIN_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_ICE_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_ICE_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_ICLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_ICLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE ICE_delayed	: STD_ULOGIC := 'X';
	VARIABLE ICLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE YIN_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_YIN_ICLK_posedge,
	 TimingData		=> Tmkr_YIN_ICLK_posedge,
	 TestSignal		=> YIN_ipd,
	 TestSignalName		=> "YIN",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName	        => "ICLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_YIN_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_YIN_ICLK_negedge_posedge,
	 HoldHigh		=> thold_YIN_ICLK_posedge_posedge,
	 HoldLow		=> thold_YIN_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (ICE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOIN_IREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_ICE_ICLK_posedge,
	 TimingData		=> Tmkr_ICE_ICLK_posedge,
	 TestSignal		=> ICE_ipd,
	 TestSignalName		=> "ICE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName		=> "ICLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_ICE_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_ICE_ICLK_negedge_posedge,
	 HoldHigh		=> thold_ICE_ICLK_posedge_posedge,
	 HoldLow		=> thold_ICE_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_ICLK_posedge,
	 TimingData		=> Tmkr_PRE_ICLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName		=> "ICLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_ICLK_negedge_posedge,
	 Removal		=> thold_PRE_ICLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((ICE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_ICLK,
	 PeriodData		=> PInfo_ICLK,
	 TestSignal		=> ICLK_ipd,
	 TestSignalName		=> "ICLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_ICLK_posedge,
	 PulseWidthLow		=> tpw_ICLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOIN_IREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "IOIN_IREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_YIN_ICLK_posedge or 
	 Tviol_ICE_ICLK_posedge or 
	 Tviol_PRE_ICLK_posedge or Tviol_PRE_ICLK_posedge or Pviol_PRE or Pviol_ICLK;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Y,
	 GlitchData => Y_GlitchData,
	 OutSignalName => "Y",
	 OutTemp => Y_zd,
	 Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_Y, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOIN_IREP_VITAL of IOIN_IREP is
   for VITAL_ACT
   end for;
end CFG_IOIN_IREP_VITAL;



 ---- CELL IOTRI_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_EB is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_DOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		DOUT		: out    STD_ULOGIC;
		EOUT		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_OB_EB :  entity is TRUE;
 end IOTRI_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        DOUT_zd :=TO_X01(D_ipd);
        EOUT_zd :=TO_X01(E_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => DOUT,
	   GlitchData => DOUT_GlitchData,
	   OutSignalName => "DOUT",
	   OutTemp => DOUT_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_DOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => EOUT,
	   GlitchData => EOUT_GlitchData,
	   OutSignalName => "EOUT",
	   OutTemp => EOUT_zd,
	   Paths => (
	             0 => (E_ipd'last_event,tpd_E_EOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOTRI_OB_EB_VITAL of IOTRI_OB_EB is 
    for VITAL_ACT
    end for;
 end CFG_IOTRI_OB_EB_VITAL;



 ---- CELL IOTRI_OB_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_ERC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OB_ERC :  entity is TRUE;
 end IOTRI_OB_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_ERC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, CLR_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_E_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS EOUT_zd : STD_LOGIC is Results(1);
	ALIAS DOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_OCLK_posedge,
	 TimingData		=> Tmkr_E_OCLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_E_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_E_OCLK_negedge_posedge,
	 HoldHigh		=> thold_E_OCLK_posedge_posedge,
	 HoldLow		=> thold_E_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OB_ERC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_OCLK_posedge,
	 TimingData             => Tmkr_CLR_OCLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => OCLK_ipd,
	 RefSignalName          => "OCLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_OCLK_negedge_posedge,
	 Removal               => thold_CLR_OCLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOTRI_OB_ERC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_E_OCLK_posedge or 
	 Pviol_CLR or 
	 Pviol_OCLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
    --- combinatorial output logic. 
   DOUT_zd :=  TO_X01(D_ipd) ;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (
	         0 => (D_ipd'last_event, tpd_D_DOUT, true),
		 1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OB_ERC_VITAL of IOTRI_OB_ERC is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OB_ERC_VITAL;



 ---- CELL IOTRI_OB_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_ERP is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OB_ERP :  entity is TRUE;
 end IOTRI_OB_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_ERP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, PRE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_E_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS EOUT_zd : STD_LOGIC is Results(1);
	ALIAS DOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_OCLK_posedge,
	 TimingData		=> Tmkr_E_OCLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_E_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_E_OCLK_negedge_posedge,
	 HoldHigh		=> thold_E_OCLK_posedge_posedge,
	 HoldLow		=> thold_E_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OB_ERP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_OCLK_posedge,
	 TimingData		=> Tmkr_PRE_OCLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_OCLK_negedge_posedge,
	 Removal		=> thold_PRE_OCLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_E_OCLK_posedge or 
	 Tviol_PRE_OCLK_posedge or 
	 Tviol_PRE_OCLK_posedge or Pviol_PRE or Pviol_OCLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
    --- combinatorial output logic. 
   DOUT_zd := TO_X01(D_ipd) ;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (
	         0 => (D_ipd'last_event, tpd_D_DOUT, true),
		 1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OB_ERP_VITAL of IOTRI_OB_ERP is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OB_ERP_VITAL;



 ---- CELL IOTRI_OB_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_EREC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OB_EREC :  entity is TRUE;
 end IOTRI_OB_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_EREC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (OCE_ipd,OCE, tipd_OCE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, CLR_ipd,OCE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_E_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_OCE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_OCE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCE_delayed	: STD_ULOGIC := 'X';
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS EOUT_zd : STD_LOGIC is Results(1);
	ALIAS DOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_OCLK_posedge,
	 TimingData		=> Tmkr_E_OCLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_E_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_E_OCLK_negedge_posedge,
	 HoldHigh		=> thold_E_OCLK_posedge_posedge,
	 HoldLow		=> thold_E_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (OCE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OB_EREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_OCE_OCLK_posedge,
	 TimingData		=> Tmkr_OCE_OCLK_posedge,
	 TestSignal		=> OCE_ipd,
	 TestSignalName		=> "OCE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_OCE_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_OCE_OCLK_negedge_posedge,
	 HoldHigh		=> thold_OCE_OCLK_posedge_posedge,
	 HoldLow		=> thold_OCE_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_OCLK_posedge,
	 TimingData             => Tmkr_CLR_OCLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => OCLK_ipd,
	 RefSignalName          => "OCLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_OCLK_negedge_posedge,
	 Removal               => thold_CLR_OCLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((OCE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOTRI_OB_EREC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_E_OCLK_posedge or 
	 Tviol_OCE_OCLK_posedge or 
	 Pviol_CLR or Pviol_OCLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
    --- combinatorial output logic. 
   DOUT_zd := TO_X01( D_ipd) ;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (
	         0 => (D_ipd'last_event, tpd_D_DOUT, true),
		 1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OB_EREC_VITAL of IOTRI_OB_EREC is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OB_EREC_VITAL;



 ---- CELL IOTRI_OB_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_EREP is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OB_EREP :  entity is TRUE;
 end IOTRI_OB_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_EREP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (OCE_ipd,OCE, tipd_OCE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, PRE_ipd,OCE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_E_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_OCE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_OCE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCE_delayed	: STD_ULOGIC := 'X';
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS EOUT_zd : STD_LOGIC is Results(1);
	ALIAS DOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_OCLK_posedge,
	 TimingData		=> Tmkr_E_OCLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_E_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_E_OCLK_negedge_posedge,
	 HoldHigh		=> thold_E_OCLK_posedge_posedge,
	 HoldLow		=> thold_E_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (OCE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OB_EREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_OCE_OCLK_posedge,
	 TimingData		=> Tmkr_OCE_OCLK_posedge,
	 TestSignal		=> OCE_ipd,
	 TestSignalName		=> "OCE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_OCE_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_OCE_OCLK_negedge_posedge,
	 HoldHigh		=> thold_OCE_OCLK_posedge_posedge,
	 HoldLow		=> thold_OCE_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_OCLK_posedge,
	 TimingData		=> Tmkr_PRE_OCLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_OCLK_negedge_posedge,
	 Removal		=> thold_PRE_OCLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((OCE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_OB_EREP",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_E_OCLK_posedge or 
	 Tviol_OCE_OCLK_posedge or 
	 Tviol_PRE_OCLK_posedge or Tviol_PRE_OCLK_posedge or Pviol_PRE or Pviol_OCLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
    --- combinatorial output logic. 
   DOUT_zd := TO_X01( D_ipd) ;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (
	         0 => (D_ipd'last_event, tpd_D_DOUT, true),
		 1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OB_EREP_VITAL of IOTRI_OB_EREP is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OB_EREP_VITAL;



 ---- CELL IOTRI_ORC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_ORC_EB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_ORC_EB :  entity is TRUE;
 end IOTRI_ORC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_ORC_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLR_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_OCLK_posedge,
	 TimingData		=> Tmkr_D_OCLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_D_OCLK_negedge_posedge,
	 HoldHigh		=> thold_D_OCLK_posedge_posedge,
	 HoldLow		=> thold_D_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_ORC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_OCLK_posedge,
	 TimingData             => Tmkr_CLR_OCLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => OCLK_ipd,
	 RefSignalName          => "OCLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_OCLK_negedge_posedge,
	 Removal               => thold_CLR_OCLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_ORC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_ORC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOTRI_ORC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_OCLK_posedge or 
	 Pviol_CLR or 
	 Pviol_OCLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
    --- combinatorial output logic. 
   EOUT_zd := TO_X01(E_ipd) ;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (
	         0 => (E_ipd'last_event, tpd_E_EOUT, true),
		 1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_ORC_EB_VITAL of IOTRI_ORC_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_ORC_EB_VITAL;



 ---- CELL IOTRI_ORP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_ORP_EB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_ORP_EB :  entity is TRUE;
 end IOTRI_ORP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_ORP_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PRE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_OCLK_posedge,
	 TimingData		=> Tmkr_D_OCLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_D_OCLK_negedge_posedge,
	 HoldHigh		=> thold_D_OCLK_posedge_posedge,
	 HoldLow		=> thold_D_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_ORP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_OCLK_posedge,
	 TimingData		=> Tmkr_PRE_OCLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_OCLK_negedge_posedge,
	 Removal		=> thold_PRE_OCLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TRUE,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_ORP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_ORP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_ORP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_OCLK_posedge or 
	 Tviol_PRE_OCLK_posedge or 
	 Tviol_PRE_OCLK_posedge or Pviol_PRE or Pviol_OCLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
    --- combinatorial output logic. 
   EOUT_zd :=  TO_X01(E_ipd) ;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (
	         0 => (E_ipd'last_event, tpd_E_EOUT, true),
		 1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_ORP_EB_VITAL of IOTRI_ORP_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_ORP_EB_VITAL;



 ---- CELL IOTRI_OREC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OREC_EB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OREC_EB :  entity is TRUE;
 end IOTRI_OREC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OREC_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (OCE_ipd,OCE, tipd_OCE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLR_ipd,OCE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_OCE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_OCE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCE_delayed	: STD_ULOGIC := 'X';
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_OCLK_posedge,
	 TimingData		=> Tmkr_D_OCLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_D_OCLK_negedge_posedge,
	 HoldHigh		=> thold_D_OCLK_posedge_posedge,
	 HoldLow		=> thold_D_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (OCE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OREC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_OCE_OCLK_posedge,
	 TimingData		=> Tmkr_OCE_OCLK_posedge,
	 TestSignal		=> OCE_ipd,
	 TestSignalName		=> "OCE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_OCE_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_OCE_OCLK_negedge_posedge,
	 HoldHigh		=> thold_OCE_OCLK_posedge_posedge,
	 HoldLow		=> thold_OCE_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT CLR_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OREC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_OCLK_posedge,
	 TimingData             => Tmkr_CLR_OCLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => OCLK_ipd,
	 RefSignalName          => "OCLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_OCLK_negedge_posedge,
	 Removal               => thold_CLR_OCLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01((OCE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OREC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_OREC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => TRUE,
	 HeaderMsg              => InstancePath & "IOTRI_OREC_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_OCLK_posedge or 
	 Tviol_OCE_OCLK_posedge or 
	 Pviol_CLR or Pviol_OCLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
    --- combinatorial output logic. 
   EOUT_zd := TO_X01(E_ipd) ;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (
	         0 => (E_ipd'last_event, tpd_E_EOUT, true),
		 1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OREC_EB_VITAL of IOTRI_OREC_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OREC_EB_VITAL;



 ---- CELL IOTRI_OREP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OREP_EB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_PRE_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_PRE_posedge		:  VitalDelayType := 0.000 ns;
		tipd_PRE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PRE		:   in    STD_ULOGIC;
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OREP_EB :  entity is TRUE;
 end IOTRI_OREP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OREP_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (PRE_ipd,PRE, tipd_PRE);
	  VitalWireDelay (OCE_ipd,OCE, tipd_OCE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PRE_ipd,OCE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_OCE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_OCE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_PRE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_PRE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
	VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCE_delayed	: STD_ULOGIC := 'X';
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_OCLK_posedge,
	 TimingData		=> Tmkr_D_OCLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_D_OCLK_negedge_posedge,
	 HoldHigh		=> thold_D_OCLK_posedge_posedge,
	 HoldLow		=> thold_D_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT PRE_ipd) AND (OCE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OREP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_OCE_OCLK_posedge,
	 TimingData		=> Tmkr_OCE_OCLK_posedge,
	 TestSignal		=> OCE_ipd,
	 TestSignalName		=> "OCE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_OCE_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_OCE_OCLK_negedge_posedge,
	 HoldHigh		=> thold_OCE_OCLK_posedge_posedge,
	 HoldLow		=> thold_OCE_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01((( NOT PRE_ipd)) ) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OREP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_PRE_OCLK_posedge,
	 TimingData		=> Tmkr_PRE_OCLK_posedge,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_PRE_OCLK_negedge_posedge,
	 Removal		=> thold_PRE_OCLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01((OCE_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OREP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT PRE_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "IOTRI_OREP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_PRE,
	 PeriodData		=> PInfo_PRE,
	 TestSignal		=> PRE_ipd,
	 TestSignalName		=> "PRE",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_PRE_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_OREP_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_OCLK_posedge or 
	 Tviol_OCE_OCLK_posedge or 
	 Tviol_PRE_OCLK_posedge or Tviol_PRE_OCLK_posedge or Pviol_PRE or Pviol_OCLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
    --- combinatorial output logic. 
   EOUT_zd := TO_X01(E_ipd) ;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
	             1=> (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (
	         0 => (E_ipd'last_event, tpd_E_EOUT, true),
		 1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true),
	           2 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OREP_EB_VITAL of IOTRI_OREP_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OREP_EB_VITAL;



 ---- CELL IOTRI_ORC_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_ORC_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_ORC_ERC :  entity is TRUE;
 end IOTRI_ORC_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_ORC_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, E_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOTRI_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOTRI_ORC_ERC_VITAL of IOTRI_ORC_ERC is
   for VITAL_ACT
   end for;
end CFG_IOTRI_ORC_ERC_VITAL;



 ---- CELL IOTRI_OREC_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OREC_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_OREC_EREC :  entity is TRUE;
 end IOTRI_OREC_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OREC_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, E_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOTRI_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OREC_EREC_VITAL of IOTRI_OREC_EREC is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OREC_EREC_VITAL;



 ---- CELL IOTRI_ORP_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_ORP_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_ORP_ERP :  entity is TRUE;
 end IOTRI_ORP_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_ORP_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, PRE_ipd, E_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOTRI_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOTRI_ORP_ERP_VITAL of IOTRI_ORP_ERP is
   for VITAL_ACT
   end for;
end CFG_IOTRI_ORP_ERP_VITAL;



 ---- CELL IOTRI_OREP_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OREP_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_OREP_EREP :  entity is TRUE;
 end IOTRI_OREP_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OREP_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, E_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow               => TRUE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOTRI_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OREP_EREP_VITAL of IOTRI_OREP_EREP is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OREP_EREP_VITAL;



 ---- CELL IOBI_IB_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_EB is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_D_DOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		YIN		: in    STD_ULOGIC;
		DOUT		: out    STD_ULOGIC;
		EOUT		: out    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_EB :  entity is TRUE;
 end IOBI_IB_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, YIN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);
	ALIAS Y_zd : STD_LOGIC is Results(3);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        DOUT_zd :=TO_X01(D_ipd);
        EOUT_zd :=TO_X01(E_ipd);
        Y_zd :=TO_X01(YIN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => DOUT,
	   GlitchData => DOUT_GlitchData,
	   OutSignalName => "DOUT",
	   OutTemp => DOUT_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_DOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => EOUT,
	   GlitchData => EOUT_GlitchData,
	   OutSignalName => "EOUT",
	   OutTemp => EOUT_zd,
	   Paths => (
	             0 => (E_ipd'last_event,tpd_E_EOUT, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (YIN_ipd'last_event,tpd_YIN_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBI_IB_OB_EB_VITAL of IOBI_IB_OB_EB is 
    for VITAL_ACT
    end for;
 end CFG_IOBI_IB_OB_EB_VITAL;



 ---- CELL IOBI_IB_OB_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_ERC :  entity is TRUE;
 end IOBI_IB_OB_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, CLR_ipd, YIN_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow               =>FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

   Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OB_ERC_VITAL of IOBI_IB_OB_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OB_ERC_VITAL;



 ---- CELL IOBI_IB_OB_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_EREC :  entity is TRUE;
 end IOBI_IB_OB_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, YIN_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OB_EREC_VITAL of IOBI_IB_OB_EREC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OB_EREC_VITAL;



 ---- CELL IOBI_IB_OB_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_ERP :  entity is TRUE;
 end IOBI_IB_OB_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, PRE_ipd, YIN_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Pviol_PRE;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OB_ERP_VITAL of IOBI_IB_OB_ERP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OB_ERP_VITAL;



 ---- CELL IOBI_IB_OB_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_EREP :  entity is TRUE;
 end IOBI_IB_OB_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, YIN_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Pviol_PRE;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OB_EREP_VITAL of IOBI_IB_OB_EREP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OB_EREP_VITAL;


---- CELL IOBI_IB_OD_EB ----
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
 entity IOBI_IB_OD_EB is
   generic (
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;

      tipd_DR          : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DF          : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E           : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_OCLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_YIN         : VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_E_EOUT       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_YIN_Y        : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLR_DOUT     : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_OCLK_DOUT    : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_DR_OCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DR_OCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_DR_OCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DR_OCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

      tsetup_DF_OCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DF_OCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_DF_OCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_DF_OCLK_negedge_posedge      : VitalDelayType := 0.000 ns;

      trecovery_CLR_OCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_CLR_OCLK_negedge_posedge     : VitalDelayType := 0.000 ns;

      tpw_OCLK_posedge                   :  VitalDelayType := 0.000 ns;
      tpw_OCLK_negedge                   :  VitalDelayType := 0.000 ns;
      tperiod_OCLK_posedge               :  VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                    :  VitalDelayType := 0.000 ns
     );


   port (
      DR            :  in    std_ulogic;
      DF            :  in    std_ulogic;
      CLR           :  in    std_ulogic;
      E             :  in    std_ulogic;
      OCLK          :  in    std_ulogic;
      YIN           :  in    std_ulogic;
      DOUT          :  out   std_ulogic;
      EOUT          :  out   std_ulogic;
      Y             :  out   std_ulogic
     );

   attribute VITAL_LEVEL0 of IOBI_IB_OD_EB :  entity is TRUE;
   
end IOBI_IB_OD_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OD_EB is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

  signal DR_ipd   : std_ulogic := 'X';
  signal DF_ipd   : std_ulogic := 'X';
  signal CLR_ipd  : std_ulogic := 'X';
  signal E_ipd    : std_ulogic := 'X';
  signal OCLK_ipd : std_ulogic := 'X';
  signal YIN_ipd  : std_ulogic := 'X';

  begin  --  VITAL_ACT
  
  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WireDelay: block

  begin  --  block WireDelay
  
    VitalWireDelay (DR_ipd,   DR,   VitalExtendToFillDelay(tipd_DR));
    VitalWireDelay (DF_ipd,   DF,   VitalExtendToFillDelay(tipd_DF));
    VitalWireDelay (CLR_ipd,  CLR,  VitalExtendToFillDelay(tipd_CLR));
    VitalWireDelay (E_ipd,    E,    VitalExtendToFillDelay(tipd_E));
    VitalWireDelay (OCLK_ipd, OCLK, VitalExtendToFillDelay(tipd_OCLK));
    VitalWireDelay (YIN_ipd,  YIN,  VitalExtendToFillDelay(tipd_YIN));

  end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################
  VITALBehavior : process (DR_ipd, DF_ipd, CLR_ipd, E_ipd, OCLK_ipd, YIN_ipd)


    -- timing check results
    variable Tviol_DR_OCLK_posedge  : std_ulogic := '0';
    variable Tmkr_DR_OCLK_posedge   : VitalTimingDataType := VitalTimingDataInit;
    variable Tviol_DF_OCLK_posedge  : std_ulogic := '0';
    variable Tmkr_DF_OCLK_posedge   : VitalTimingDataType := VitalTimingDataInit;
    variable Tviol_CLR_OCLK_posedge : std_ulogic := '0';
    variable Tmkr_CLR_OCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
    variable Pviol_OCLK             : std_ulogic := '0';
    variable PInfo_OCLK             : VitalPeriodDataType := VitalPeriodDataInit;
    variable Pviol_CLR              : std_ulogic := '0';
    variable PInfo_CLR              : VitalPeriodDataType := VitalPeriodDataInit;

    -- functionality results
    variable Violation              : std_ulogic := '0';
    variable PrevData_DR            : STD_LOGIC_VECTOR(0 to 2);
    variable PrevData_DF            : STD_LOGIC_VECTOR(0 to 2);

    variable DOUT_zd                : std_ulogic := 'X';
    variable EOUT_zd                : std_ulogic := 'X';
    variable tmp1_zd                : std_ulogic := 'X';
    variable tmp2_zd                : std_ulogic := 'X';
    variable Y_zd                   : std_ulogic := 'X';

    -- output glitch detection variables
    variable DOUT_GlitchData        : VitalGlitchDataType;
    variable EOUT_GlitchData        : VitalGlitchDataType;
    variable Y_GlitchData           : VitalGlitchDataType;

  begin
  
    ------------------------
    --  Timing Check Section
    ------------------------

    if (TimingChecksOn) then
       VitalSetupHoldCheck (
         Violation              => Tviol_DR_OCLK_posedge,
         TimingData             => Tmkr_DR_OCLK_posedge,
         TestSignal             => DR_ipd,
         TestSignalName         => "DR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DR_OCLK_posedge_posedge,
         SetupLow               => tsetup_DR_OCLK_negedge_posedge,
         HoldHigh               => thold_DR_OCLK_posedge_posedge,
         HoldLow                => thold_DR_OCLK_negedge_posedge,
         CheckEnabled           => TO_X01(CLR_ipd) /= '1',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_IB_OD_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_DF_OCLK_posedge,
         TimingData             => Tmkr_DF_OCLK_posedge,
         TestSignal             => DF_ipd,
         TestSignalName         => "DF",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DF_OCLK_posedge_posedge,
         SetupLow               => tsetup_DF_OCLK_negedge_posedge,
         HoldHigh               => thold_DF_OCLK_posedge_posedge,
         HoldLow                => thold_DF_OCLK_negedge_posedge,
         CheckEnabled           => TO_X01(CLR_ipd) /= '1',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_IB_OD_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

       VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_OCLK_posedge,
         TimingData             => Tmkr_CLR_OCLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         Recovery               => trecovery_CLR_OCLK_negedge_posedge,
         Removal                => thold_CLR_OCLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_IB_OD_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

       VitalPeriodPulseCheck (
         Violation              => Pviol_OCLK,
         PeriodData             => PInfo_OCLK,
         TestSignal             => OCLK_ipd,
         TestSignalName         => "OCLK",
         TestDelay              => 0 ns,
         Period                 => tperiod_OCLK_posedge,
         PulseWidthHigh         => tpw_OCLK_posedge,
         PulseWidthLow          => tpw_OCLK_negedge,
         CheckEnabled           => TO_X01(CLR_ipd) /= '1',
         HeaderMsg              => InstancePath & "/IOBI_IB_OD_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);


       VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period                 => 0 ns,
         PulseWidthHigh         => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOBI_IB_OD_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

    end if;
    
    --------------------------------
    --  Functionality Section
    -------------------------------

    Violation := Tviol_DR_OCLK_posedge or Tviol_DF_OCLK_posedge or 
                 Tviol_CLR_OCLK_posedge or Pviol_OCLK or Pviol_CLR;

    Y_zd    := TO_X01(YIN_ipd);
    EOUT_zd := TO_X01(E_ipd);

    VitalStateTable(
      Result => tmp1_zd,
      PreviousDataIn => PrevData_DR,
      StateTable => DFN1C1_Q_tab,
      DataIn => ( CLR_ipd, OCLK_ipd, DR_ipd ));
    tmp1_zd := Violation XOR tmp1_zd;

    VitalStateTable(
      Result => tmp2_zd,
      PreviousDataIn => PrevData_DF,
      StateTable => DFN1C1_Q_tab,
      DataIn => ( CLR_ipd, OCLK_ipd, DF_ipd ));
    tmp2_zd := Violation XOR tmp2_zd;

    DOUT_zd := VitalMUX2(tmp1_zd, tmp2_zd, OCLK_ipd);

    ----------------------
    --  Path Delay Section
    ----------------------
    
    VitalPathDelay01 (
         OutSignal     => DOUT,
         GlitchData    => DOUT_GlitchData,
         OutSignalName => "DOUT",
         OutTemp       => DOUT_zd,
         Paths         => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
                           1 => (CLR_ipd'last_event,  tpd_CLR_DOUT,  true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

    VitalPathDelay01 (
         OutSignal     => EOUT,
         GlitchData    => EOUT_GlitchData,
         OutSignalName => "EOUT",
         OutTemp       => EOUT_zd,
         Paths         => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

    VitalPathDelay01 (
         OutSignal     => Y,
         GlitchData    => Y_GlitchData,
         OutSignalName => "Y",
         OutTemp       => Y_zd,
         Paths         => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

  end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OD_EB_VITAL of IOBI_IB_OD_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OD_EB_VITAL;

 ---- CELL IOBI_IB_ORC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_ORC_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_ORC_EB :  entity is TRUE;
 end IOBI_IB_ORC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_ORC_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, CLR_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_ORC_EB_VITAL of IOBI_IB_ORC_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_ORC_EB_VITAL;



 ---- CELL IOBI_IB_OREC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OREC_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OREC_EB :  entity is TRUE;
 end IOBI_IB_OREC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OREC_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OREC_EB_VITAL of IOBI_IB_OREC_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OREC_EB_VITAL;



 ---- CELL IOBI_IB_ORP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_ORP_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_ORP_EB :  entity is TRUE;
 end IOBI_IB_ORP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_ORP_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, PRE_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Pviol_PRE;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_ORP_EB_VITAL of IOBI_IB_ORP_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_ORP_EB_VITAL;



 ---- CELL IOBI_IB_OREP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OREP_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OREP_EB :  entity is TRUE;
 end IOBI_IB_OREP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OREP_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Pviol_PRE;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OREP_EB_VITAL of IOBI_IB_OREP_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OREP_EB_VITAL;



 ---- CELL IOBI_IB_ORC_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_ORC_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_ORC_ERC :  entity is TRUE;
 end IOBI_IB_ORC_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_ORC_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, E_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_ORC_ERC_VITAL of IOBI_IB_ORC_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_ORC_ERC_VITAL;



 ---- CELL IOBI_IB_OREC_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OREC_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OREC_EREC :  entity is TRUE;
 end IOBI_IB_OREC_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OREC_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, E_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OREC_EREC_VITAL of IOBI_IB_OREC_EREC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OREC_EREC_VITAL;



 ---- CELL IOBI_IB_ORP_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_ORP_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_ORP_ERP :  entity is TRUE;
 end IOBI_IB_ORP_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_ORP_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, PRE_ipd, E_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_ORP_ERP_VITAL of IOBI_IB_ORP_ERP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_ORP_ERP_VITAL;



 ---- CELL IOBI_IB_OREP_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OREP_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OREP_EREP :  entity is TRUE;
 end IOBI_IB_OREP_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OREP_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, E_ipd, YIN_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IB_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

        Y_zd :=TO_X01(YIN_ipd);


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OREP_EREP_VITAL of IOBI_IB_OREP_EREP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OREP_EREP_VITAL;



 ---- CELL IOBI_IRC_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_OB_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_OB_EB :  entity is TRUE;
 end IOBI_IRC_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_OB_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, YIN_ipd, ICLK_ipd, CLR_ipd)


   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_CLR_ICLK_posedge  or Pviol_CLR;

        DOUT_zd :=TO_X01(D_ipd);

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_OB_EB_VITAL of IOBI_IRC_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_OB_EB_VITAL;



 ---- CELL IOBI_IREC_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_OB_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_OB_EB :  entity is TRUE;
 end IOBI_IREC_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_OB_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, YIN_ipd, ICLK_ipd, CLR_ipd, ICE_ipd)


   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_OB_EB_VITAL of IOBI_IREC_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_OB_EB_VITAL;



 ---- CELL IOBI_IRP_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_OB_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_OB_EB :  entity is TRUE;
 end IOBI_IRP_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_OB_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, YIN_ipd, ICLK_ipd, PRE_ipd)


   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_PRE_ICLK_posedge  or Pviol_PRE;

        DOUT_zd :=TO_X01(D_ipd);

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_OB_EB_VITAL of IOBI_IRP_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_OB_EB_VITAL;



 ---- CELL IOBI_IREP_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_OB_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_OB_EB :  entity is TRUE;
 end IOBI_IREP_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_OB_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, YIN_ipd, ICLK_ipd, ICE_ipd, PRE_ipd)


   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE;

        DOUT_zd :=TO_X01(D_ipd);

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_OB_EB_VITAL of IOBI_IREP_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_OB_EB_VITAL;



 ---- CELL IOBI_IRC_OB_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_OB_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_OB_ERC :  entity is TRUE;
 end IOBI_IRC_OB_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_OB_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, CLR_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh               => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period                 => 0 ns,
    PulseWidthHigh         => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge, 
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period                 => 0 ns,
    PulseWidthHigh         => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh               => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period                 => 0 ns,
    PulseWidthHigh         => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_OB_ERC_VITAL of IOBI_IRC_OB_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_OB_ERC_VITAL;



 ---- CELL IOBI_IREC_OB_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_OB_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_OB_ERC :  entity is TRUE;
 end IOBI_IREC_OB_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_OB_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, CLR_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_OB_ERC_VITAL of IOBI_IREC_OB_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_OB_ERC_VITAL;



 ---- CELL IOBI_IRC_OB_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_OB_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_OB_EREC :  entity is TRUE;
 end IOBI_IRC_OB_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_OB_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_OB_EREC_VITAL of IOBI_IRC_OB_EREC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_OB_EREC_VITAL;



 ---- CELL IOBI_IREC_OB_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_OB_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_OB_EREC :  entity is TRUE;
 end IOBI_IREC_OB_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_OB_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OB_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OB_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_OB_EREC_VITAL of IOBI_IREC_OB_EREC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_OB_EREC_VITAL;



 ---- CELL IOBI_IRP_OB_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_OB_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_OB_ERP :  entity is TRUE;
 end IOBI_IRP_OB_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_OB_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, PRE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_OB_ERP_VITAL of IOBI_IRP_OB_ERP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_OB_ERP_VITAL;



 ---- CELL IOBI_IREP_OB_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_OB_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_OB_ERP :  entity is TRUE;
 end IOBI_IREP_OB_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_OB_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, PRE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_OB_ERP_VITAL of IOBI_IREP_OB_ERP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_OB_ERP_VITAL;



 ---- CELL IOBI_IRP_OB_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_OB_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_OB_EREP :  entity is TRUE;
 end IOBI_IRP_OB_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_OB_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_OB_EREP_VITAL of IOBI_IRP_OB_EREP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_OB_EREP_VITAL;



 ---- CELL IOBI_IREP_OB_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_OB_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_OB_EREP :  entity is TRUE;
 end IOBI_IREP_OB_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_OB_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OB_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OB_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_OB_EREP_VITAL of IOBI_IREP_OB_EREP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_OB_EREP_VITAL;



 ---- CELL IOBI_IRC_ORC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_ORC_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_ORC_EB :  entity is TRUE;
 end IOBI_IRC_ORC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_ORC_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, CLR_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);

   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_ORC_EB_VITAL of IOBI_IRC_ORC_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_ORC_EB_VITAL;



 ---- CELL IOBI_IREC_ORC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_ORC_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_ORC_EB :  entity is TRUE;
 end IOBI_IREC_ORC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_ORC_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, CLR_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);

   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_ORC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_ORC_EB_VITAL of IOBI_IREC_ORC_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_ORC_EB_VITAL;



 ---- CELL IOBI_IRC_OREC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_OREC_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_OREC_EB :  entity is TRUE;
 end IOBI_IRC_OREC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_OREC_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_OREC_EB_VITAL of IOBI_IRC_OREC_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_OREC_EB_VITAL;



 ---- CELL IOBI_IREC_OREC_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_OREC_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_OREC_EB :  entity is TRUE;
 end IOBI_IREC_OREC_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_OREC_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_OREC_EB_VITAL of IOBI_IREC_OREC_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_OREC_EB_VITAL;



 ---- CELL IOBI_IRP_ORP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_ORP_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_ORP_EB :  entity is TRUE;
 end IOBI_IRP_ORP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_ORP_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, PRE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_ORP_EB_VITAL of IOBI_IRP_ORP_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_ORP_EB_VITAL;



 ---- CELL IOBI_IRP_OREP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_OREP_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_OREP_EB :  entity is TRUE;
 end IOBI_IRP_OREP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_OREP_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_OREP_EB_VITAL of IOBI_IRP_OREP_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_OREP_EB_VITAL;



 ---- CELL IOBI_IREP_ORP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_ORP_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_ORP_EB :  entity is TRUE;
 end IOBI_IREP_ORP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_ORP_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, PRE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_ORP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_ORP_EB_VITAL of IOBI_IREP_ORP_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_ORP_EB_VITAL;



 ---- CELL IOBI_IREP_OREP_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_OREP_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_OREP_EB :  entity is TRUE;
 end IOBI_IREP_OREP_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_OREP_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_OREP_EB_VITAL of IOBI_IREP_OREP_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_OREP_EB_VITAL;



 ---- CELL IOBI_IRC_ORC_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_ORC_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_ORC_ERC :  entity is TRUE;
 end IOBI_IRC_ORC_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_ORC_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, E_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_ORC_ERC_VITAL of IOBI_IRC_ORC_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_ORC_ERC_VITAL;



 ---- CELL IOBI_IRC_OREC_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRC_OREC_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRC_OREC_EREC :  entity is TRUE;
 end IOBI_IRC_OREC_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRC_OREC_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, E_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRC_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRC_OREC_EREC_VITAL of IOBI_IRC_OREC_EREC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRC_OREC_EREC_VITAL;



 ---- CELL IOBI_IREC_ORC_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_ORC_ERC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_ORC_ERC :  entity is TRUE;
 end IOBI_IREC_ORC_ERC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_ORC_ERC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, E_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_ORC_ERC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_ORC_ERC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_ORC_ERC_VITAL of IOBI_IREC_ORC_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_ORC_ERC_VITAL;



 ---- CELL IOBI_IREC_OREC_EREC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREC_OREC_EREC is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_CLR_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_CLR_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                CLR         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREC_OREC_EREC :  entity is TRUE;
 end IOBI_IREC_OREC_EREC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREC_OREC_EREC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, CLR_ipd, OCE_ipd, E_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLR    : STD_ULOGIC := '0';
   VARIABLE PInfo_CLR    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE CLR_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_OCLK_posedge,
   TimingData             => Tmkr_CLR_OCLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_OCLK_negedge_posedge,
   Removal                => thold_CLR_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_CLR,
    PeriodData             => PInfo_CLR,
    TestSignal             => CLR_ipd,
    TestSignalName         => "CLR",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_CLR_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_CLR_ICLK_posedge,
   TimingData             => Tmkr_CLR_ICLK_posedge,
   TestSignal             => CLR_ipd,
   TestSignalName         => "CLR",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_CLR_ICLK_negedge_posedge,
   Removal                => thold_CLR_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREC_OREC_EREC",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREC_OREC_EREC",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_CLR_OCLK_posedge  or Tviol_CLR_ICLK_posedge  or Pviol_CLR or Tviol_OCE_OCLK_posedge  or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (CLR_ipd'last_event, tpd_CLR_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREC_OREC_EREC_VITAL of IOBI_IREC_OREC_EREC is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREC_OREC_EREC_VITAL;



 ---- CELL IOBI_IRP_ORP_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_ORP_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_ORP_ERP :  entity is TRUE;
 end IOBI_IRP_ORP_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_ORP_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, PRE_ipd, E_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_ORP_ERP_VITAL of IOBI_IRP_ORP_ERP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_ORP_ERP_VITAL;



 ---- CELL IOBI_IRP_OREP_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRP_OREP_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRP_OREP_EREP :  entity is TRUE;
 end IOBI_IRP_OREP_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRP_OREP_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, E_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRP_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRP_OREP_EREP_VITAL of IOBI_IRP_OREP_EREP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRP_OREP_EREP_VITAL;



 ---- CELL IOBI_IREP_ORP_ERP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_ORP_ERP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_ORP_ERP :  entity is TRUE;
 end IOBI_IREP_ORP_ERP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_ORP_ERP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, PRE_ipd, E_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_ORP_ERP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_ORP_ERP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_ORP_ERP_VITAL of IOBI_IREP_ORP_ERP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_ORP_ERP_VITAL;



 ---- CELL IOBI_IREP_OREP_EREP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IREP_OREP_EREP is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PRE_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		trecovery_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_OCLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tpw_PRE_posedge	:  VitalDelayType := 0.000 ns;
		trecovery_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_PRE_ICLK_negedge_posedge	:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PRE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                PRE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IREP_OREP_EREP :  entity is TRUE;
 end IOBI_IREP_OREP_EREP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IREP_OREP_EREP is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, OCLK_ipd, OCE_ipd, PRE_ipd, E_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_PRE    : STD_ULOGIC := '0';
   VARIABLE PInfo_PRE    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q0  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE PRE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_OCLK_posedge,
   TimingData             => Tmkr_PRE_OCLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_OCLK_negedge_posedge,
   Removal                => thold_PRE_OCLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_PRE,
    PeriodData             => PInfo_PRE,
    TestSignal             => PRE_ipd,
    TestSignalName         => "PRE",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_PRE_posedge,
    PulseWidthLow          => 0 ns,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalRecoveryRemovalCheck  (
   Violation              => Tviol_PRE_ICLK_posedge,
   TimingData             => Tmkr_PRE_ICLK_posedge,
   TestSignal             => PRE_ipd,
   TestSignalName         => "PRE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   Recovery               => trecovery_PRE_ICLK_negedge_posedge,
   Removal                => thold_PRE_ICLK_negedge_posedge,
   ActiveLow              => FALSE,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IREP_OREP_EREP",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IREP_OREP_EREP",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_PRE_OCLK_posedge  or Tviol_PRE_ICLK_posedge  or Pviol_PRE or Tviol_E_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q0,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), (NOT PRE_ipd), OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), (NOT PRE_ipd), ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;
   E_delayed := E_ipd;

   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
              1 => (PRE_ipd'last_event, tpd_PRE_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true),
              1 => (PRE_ipd'last_event, tpd_PRE_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IREP_OREP_EREP_VITAL of IOBI_IREP_OREP_EREP is
   for VITAL_ACT
   end for;
end CFG_IOBI_IREP_OREP_EREP_VITAL;



 ---- CELL IOPAD_IN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_IN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_IN :  entity is TRUE;
 end IOPAD_IN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_IN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

        -- timing check results
        VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_IN_VITAL of IOPAD_IN is 
    for VITAL_ACT
    end for;

 end CFG_IOPAD_IN_VITAL;



 ---- CELL IOPADP_BI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPADP_BI is
    generic(
       TimingChecksOn : Boolean  := True;
       Xon            : Boolean  := False;
       InstancePath   : STRING   := "*";
       MsgOn          : Boolean  := True;

                tpw_D_posedge     : VitalDelayType    := 0.000 ns;
                tpw_D_negedge     : VitalDelayType    := 0.000 ns;
                tpw_E_posedge     : VitalDelayType    := 0.000 ns;
                tpw_E_negedge     : VitalDelayType    := 0.000 ns;
                tpw_PAD_negedge   : VitalDelayType    := 0.000 ns;
                tpw_PAD_posedge   : VitalDelayType    := 0.000 ns;
                tpw_N2PIN_negedge : VitalDelayType    := 0.000 ns;
                tpw_N2PIN_posedge : VitalDelayType    := 0.000 ns;

                tpd_D_PAD         : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PAD         : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_PAD_Y         : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_N2PIN_Y       : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_D_Y           : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_Y           : VitalDelayType01  := (0.100 ns, 0.100 ns);

                tipd_D            : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_E            : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PAD          : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_N2PIN        : VitalDelayType01  := (0.000 ns, 0.000 ns));


    port(
                D               : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                N2PIN           : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                Y               : out   STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPADP_BI :  entity is TRUE;
 end IOPADP_BI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of IOPADP_BI is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

        SIGNAL D_ipd     : STD_ULOGIC := 'X';
        SIGNAL E_ipd     : STD_ULOGIC := 'X';
        SIGNAL PAD_ipd   : STD_ULOGIC := 'X';
        SIGNAL N2PIN_ipd : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay ( D_ipd,     D,     tipd_D     );
        VitalWireDelay ( E_ipd,     E,     tipd_E     );
        VitalWireDelay ( PAD_ipd  , PAD,   tipd_PAD   );
        VitalWireDelay ( N2PIN_ipd, N2PIN, tipd_N2PIN );
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (D_ipd, E_ipd, PAD_ipd, N2PIN_ipd)

        -- timing check results
        VARIABLE Pviol_D         : STD_ULOGIC := '0';
        VARIABLE PeriodData_D    : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E         : STD_ULOGIC := '0';
        VARIABLE PeriodData_E    : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_N2PIN      : STD_ULOGIC := '0';
        VARIABLE PeriodData_N2PIN : VitalPeriodDataType := VitalPeriodDataInit;


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS PAD_zd     : STD_LOGIC is Results(1);
        ALIAS Y_zd       : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData  : VitalGlitchDataType;
        VARIABLE Y_GlitchData     : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_N2PIN,
              PeriodData     => PeriodData_N2PIN,
              TestSignal     => N2PIN_ipd,
              TestSignalName => "N2PIN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_N2PIN_posedge,
              PulseWidthLow  => tpw_N2PIN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


       -------------------------
       --  Functionality Section
       -------------------------
       PAD_zd   := VitalBUFIF0 (data => D_ipd, enable =>(NOT E_ipd));

       if ( TO_X01 ( PAD_ipd ) = '1' and TO_X01 ( N2PIN_ipd ) = '0' ) then
         Y_zd   := '1';
       elsif ( TO_X01 ( PAD_ipd ) = '0' and TO_X01 ( N2PIN_ipd ) = '1' ) then
         Y_zd   := '0';
       else
         Y_zd   := 'X';
       end if;


       ----------------------
       --  Path Delay Section
       ----------------------

       VitalPathDelay01Z (
         OutSignal     => PAD,
         GlitchData    => PAD_GlitchData,
         OutSignalName => "PAD",
         OutTemp       => PAD_zd,
         Paths    => (
                     0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
                     1 => (E_ipd'last_event,tpd_E_PAD, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING,
         OutputMap     => "UX01ZWLH-");

       VitalPathDelay01 (
         OutSignal     => Y,
         GlitchData    => Y_GlitchData,
         OutSignalName => "Y",
         OutTemp       => Y_zd,
         Paths    => (
                     0 => (D_ipd'last_event,tpd_D_Y, true),
                     1 => (E_ipd'last_event,tpd_E_Y, true),
                     2 => (PAD_ipd'last_event,tpd_PAD_Y, true),
                     3 => (N2PIN_ipd'last_event,tpd_N2PIN_Y, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPADP_BI_VITAL of IOPADP_BI is
    for VITAL_ACT
    end for;
 end CFG_IOPADP_BI_VITAL;


----- CELL IOPADP_IN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
 entity IOPADP_IN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
      tpw_N2PIN_posedge         : VitalDelayType := 0.000 ns;
      tpw_N2PIN_negedge         : VitalDelayType := 0.000 ns;
      tpd_PAD_Y                      :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_N2PIN_Y                    :        VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD                       :        VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_N2PIN                     :        VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :        in    STD_ULOGIC;
      N2PIN                         :        in    STD_ULOGIC;
      Y                              :        out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADP_IN : entity is FALSE;
end IOPADP_IN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IOPADP_IN is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PAD_ipd      : STD_ULOGIC := 'X';
   SIGNAL N2PIN_ipd    : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   VitalWireDelay (N2PIN_ipd, N2PIN, tipd_N2PIN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd, N2PIN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   ALIAS X_zd : STD_LOGIC is Results(2);
  
   -- timing check results
  VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
  VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;
  VARIABLE Pviol_N2PIN       : STD_ULOGIC := '0'; 
  VARIABLE PeriodData_N2PIN  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE Y_GlitchData      : VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_N2PIN,
              PeriodData     => PeriodData_N2PIN,
              TestSignal     => PAD_ipd,
              TestSignalName => "N2PIN",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_N2PIN_posedge,
              PulseWidthLow  => tpw_N2PIN_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);
      X_zd := TO_X01(N2PIN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IOPADP_IN_VITAL of IOPADP_IN is
   for VITAL_ACT
   end for;
end CFG_IOPADP_IN_VITAL;



 ---- CELL IOPADN_BI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPADN_BI is
    generic(
       TimingChecksOn : Boolean  := True;
       Xon            : Boolean  := False;
       InstancePath   : STRING   := "*";
       MsgOn          : Boolean  := True;

                tpw_DB_posedge    : VitalDelayType    := 0.000 ns;
                tpw_DB_negedge    : VitalDelayType    := 0.000 ns;
                tpw_E_posedge     : VitalDelayType    := 0.000 ns;
                tpw_E_negedge     : VitalDelayType    := 0.000 ns;
                tpw_PAD_negedge   : VitalDelayType    := 0.000 ns;
                tpw_PAD_posedge   : VitalDelayType    := 0.000 ns;

                tpd_DB_PAD        : VitalDelayType01  := (0.100 ns, 0.100 ns);
                tpd_E_PAD         : VitalDelayType01Z := (0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns, 0.100 ns);
                tpd_PAD_N2POUT    : VitalDelayType01  := (0.100 ns, 0.100 ns);

                tipd_DB           : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_E            : VitalDelayType01  := (0.000 ns, 0.000 ns);
                tipd_PAD          : VitalDelayType01  := (0.000 ns, 0.000 ns));


    port(
                DB              : in    STD_ULOGIC;
                E               : in    STD_ULOGIC;
                PAD             : inout STD_ULOGIC;
                N2POUT          : out   STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPADN_BI :  entity is TRUE;
 end IOPADN_BI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of IOPADN_BI is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

        SIGNAL DB_ipd     : STD_ULOGIC := 'X';
        SIGNAL E_ipd      : STD_ULOGIC := 'X';
        SIGNAL PAD_ipd    : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay ( DB_ipd,    DB,    tipd_DB  );
        VitalWireDelay ( E_ipd,     E,     tipd_E   );
        VitalWireDelay ( PAD_ipd  , PAD,   tipd_PAD );
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (DB_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_DB        : STD_ULOGIC := '0';
        VARIABLE PeriodData_DB   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E         : STD_ULOGIC := '0';
        VARIABLE PeriodData_E    : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
        ALIAS PAD_zd     : STD_LOGIC is Results(1);
        ALIAS N2POUT_zd  : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE PAD_GlitchData    : VitalGlitchDataType;
        VARIABLE N2POUT_GlitchData : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_DB,
              PeriodData     => PeriodData_DB,
              TestSignal     => DB_ipd,
              TestSignalName => "DB",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_DB_posedge,
              PulseWidthLow  => tpw_DB_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


       -------------------------
       --  Functionality Section
       -------------------------
       PAD_zd := VitalBUFIF0 (data => (NOT DB_ipd), enable =>(NOT E_ipd));
       N2POUT_zd := VitalBUF (data => PAD_ipd);


       ----------------------
       --  Path Delay Section
       ----------------------

       VitalPathDelay01Z (
         OutSignal     => PAD,
         GlitchData    => PAD_GlitchData,
         OutSignalName => "PAD",
         OutTemp       => PAD_zd,
         Paths    => (
                     0 => (DB_ipd'last_event,VitalExtendToFillDelay(tpd_DB_PAD),true),
                     1 => (E_ipd'last_event,tpd_E_PAD, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING,
         OutputMap     => "UX01ZWLH-");

       VitalPathDelay01 (
         OutSignal     => N2POUT,
         GlitchData    => N2POUT_GlitchData,
         OutSignalName => "N2POUT",
         OutTemp       => N2POUT_zd,
         Paths    => (
                     0 => (PAD_ipd'last_event,tpd_PAD_N2POUT, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPADN_BI_VITAL of IOPADN_BI is
    for VITAL_ACT
    end for;
 end CFG_IOPADN_BI_VITAL;



----- CELL IOPADN_IN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
 entity IOPADN_IN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
      tpw_PAD_negedge           : VitalDelayType := 0.000 ns;      
      tpd_PAD_N2POUT                 :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      N2POUT                         :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADN_IN : entity is FALSE;
end IOPADN_IN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IOPADN_IN is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS N2POUT_zd : STD_LOGIC is Results(1);

   -- timing check results
   VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
   VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE N2POUT_GlitchData	: VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_IN",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      N2POUT_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => N2POUT,
       GlitchData => N2POUT_GlitchData,
       OutSignalName => "N2POUT",
       OutTemp => N2POUT_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_N2POUT, TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IOPADN_IN_VITAL of IOPADN_IN is
   for VITAL_ACT
   end for;
end CFG_IOPADN_IN_VITAL;


 ---- CELL IOPAD_TRI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_TRI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_D_posedge 		: VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge 	 	: VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_TRI :  entity is TRUE;
 end IOPAD_TRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_TRI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_E, 
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_D, 
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_TRI_VITAL of IOPAD_TRI is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_TRI_VITAL;



----- CELL IOPADP_TRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
 entity IOPADP_TRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_E_posedge                  :  VitalDelayType := 0.000 ns;
      tpw_E_negedge		     :  VitalDelayType := 0.000 ns;
      tpw_D_posedge		     :  VitalDelayType := 0.000 ns;
      tpw_D_negedge		     :  VitalDelayType := 0.000 ns;

      tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADP_TRI : entity is FALSE;
end IOPADP_TRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IOPADP_TRI is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   
   -- timing check results
   VARIABLE Pviol_D       : STD_ULOGIC := '0'; 
   VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_E      : STD_ULOGIC := '0'; 
   VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
           
            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADP_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_IOPADP_TRI_VITAL of IOPADP_TRI is
   for VITAL_ACT
   end for;
end CFG_IOPADP_TRI_VITAL;


----- CELL IOPADN_TRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
 entity IOPADN_TRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      
      tpw_E_posedge              : VitalDelayType := 0.000 ns;    
      tpw_E_negedge		     : VitalDelayType := 0.000 ns;
      tpw_DB_posedge	     : VitalDelayType := 0.000 ns;
      tpw_DB_negedge             : VitalDelayType := 0.000 ns;
	
      tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
      tpd_DB_PAD                     :	VitalDelayType01 := (0.100 ns, 0.100 ns);
      tipd_DB                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      DB                             :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IOPADN_TRI : entity is FALSE;
end IOPADN_TRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of IOPADN_TRI is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL DB_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (DB_ipd, DB, tipd_DB);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (DB_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- timing check results
   VARIABLE Pviol_DB      : STD_ULOGIC := '0';
   VARIABLE PeriodData_DB : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_E       : STD_ULOGIC := '0';
   VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_DB,
              PeriodData     => PeriodData_DB,
              TestSignal     => DB_ipd,
              TestSignalName => "DB",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_DB_posedge,
              PulseWidthLow  => tpw_DB_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_TRI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => (NOT DB_ipd),
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (DB_ipd'last_event, VitalExtendToFillDelay(tpd_DB_PAD), TRUE)),
       Mode => VitalTransport,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_IOPADN_TRI_VITAL of IOPADN_TRI is
   for VITAL_ACT
   end for;
end CFG_IOPADN_TRI_VITAL;


 ---- CELL IOPAD_BI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_BI is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_BI :  entity is TRUE;
 end IOPAD_BI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_BI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

        -- timing check results
	VARIABLE Pviol_D	:STD_ULOGIC := '0';
        VARIABLE PeriodData_D        :VitalPeriodDataType := VitalPeriodDataInit;
 	VARIABLE Pviol_E	:STD_ULOGIC := '0';
        VARIABLE PeriodData_E        :VitalPeriodDataType := VitalPeriodDataInit;	
        VARIABLE Pviol_PAD	:STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD        :VitalPeriodDataType := VitalPeriodDataInit;     

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
         
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
 

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
          
        end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_BI_VITAL of IOPAD_BI is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_BI_VITAL;



 ---- CELL IOPAD_IN_U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_IN_U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_PAD_posedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
                tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_IN_U :  entity is TRUE;
 end IOPAD_IN_U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_IN_U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
	VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_IN_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_IN_U_VITAL of IOPAD_IN_U is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_IN_U_VITAL;



 ---- CELL IOPAD_IN_D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_IN_D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_PAD_posedge 		: VitalDelayType := 0.000 ns;
                tpw_PAD_negedge           : VitalDelayType := 0.000 ns;
                tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_IN_D :  entity is TRUE;
 end IOPAD_IN_D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_IN_D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	
        -- timing check results
	VARIABLE Pviol_PAD       : STD_ULOGIC := '0';
	VARIABLE PeriodData_PAD  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_IN_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','L'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_IN_D_VITAL of IOPAD_IN_D is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_IN_D_VITAL;



 ---- CELL IOPAD_TRI_U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_TRI_U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge 	    : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                
                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_TRI_U :  entity is TRUE;
 end IOPAD_TRI_U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_TRI_U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
        VARIABLE PeriodData_D : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
           
           VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_TRI_U_VITAL of IOPAD_TRI_U is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_TRI_U_VITAL;



 ---- CELL IOPAD_TRI_D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_TRI_D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		
                tpw_D_posedge   : VitalDelayType := 0.000 ns;
                tpw_D_negedge   : VitalDelayType := 0.000 ns;
                tpw_E_posedge   : VitalDelayType := 0.000 ns;
                tpw_E_negedge   : VitalDelayType := 0.000 ns; 

                tpd_D_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_TRI_D :  entity is TRUE;
 end IOPAD_TRI_D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_TRI_D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- timing check results
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin
          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_TRI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_TRI_D_VITAL of IOPAD_TRI_D is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_TRI_D_VITAL;



 ---- CELL IOPAD_BI_U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_BI_U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
	
		tpw_E_posedge       : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_D_posedge       : VitalDelayType := 0.000 ns;
                tpw_D_negedge 	    : VitalDelayType := 0.000 ns;
		tpw_PAD_posedge     : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge     : VitalDelayType := 0.000 ns;

             	tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		
                tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_BI_U :  entity is TRUE;
 end IOPAD_BI_U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_BI_U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- timing check results
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE PViol_PAD     : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD :VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        if ( TimingChecksOn) then
        
        
            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
            
             VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

             VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

           end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPAD_BI_U_VITAL of IOPAD_BI_U is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_BI_U_VITAL;



 ---- CELL IOPAD_BI_D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPAD_BI_D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpw_E_posedge   : VitalDelayType := 0.000 ns;
                tpw_E_negedge 	: VitalDelayType := 0.000 ns;
		tpw_D_posedge   : VitalDelayType := 0.000 ns;
                tpw_D_negedge 	: VitalDelayType := 0.000 ns;
		tpw_PAD_posedge : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge : VitalDelayType := 0.000 ns;		

                tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
	        tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
	        tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPAD_BI_D :  entity is TRUE;
 end IOPAD_BI_D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPAD_BI_D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

        -- timing check results
	VARIABLE Pviol_D       : STD_ULOGIC := '0';
	VARIABLE PeriodData_D  : VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_E       : STD_ULOGIC := '0';
	VARIABLE PeriodData_E  : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE PViol_PAD     : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD :VitalPeriodDataType := VitalPeriodDataInit;


	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin
        
        if ( TimingChecksOn ) then
        
            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
 
            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            ); 
         
            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPAD_BI_D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );
           end if;
	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

end process;

end VITAL_ACT;

 configuration CFG_IOPAD_BI_D_VITAL of IOPAD_BI_D is 
    for VITAL_ACT
    end for;
 end CFG_IOPAD_BI_D_VITAL;

 ---- CELL IOPADN_OUT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOPADN_OUT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
                tpw_DB_posedge : VitalDelayType := 0.000 ns;
                tpw_DB_negedge : VitalDelayType := 0.000 ns;
		tpd_DB_PAD     : VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_DB        : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		DB		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOPADN_OUT :  entity is TRUE;
 end IOPADN_OUT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL_ACT of IOPADN_OUT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL DB_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (DB_ipd, DB, tipd_DB);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (DB_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

        -- timing check results
        VARIABLE Pviol_DB      : STD_ULOGIC := '0';
        VARIABLE PeriodData_DB : VitalPeriodDataType := VitalPeriodDataInit;

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

          if ( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_DB,
              PeriodData     => PeriodData_DB,
              TestSignal     => DB_ipd,
              TestSignalName => "DB",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_DB_posedge,
              PulseWidthLow  => tpw_DB_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/IOPADN_OUT",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

          end if;

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd :=  (NOT DB_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (DB_ipd'last_event,tpd_DB_PAD, true)),
	  Mode => VitalTransport,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOPADN_OUT_VITAL of IOPADN_OUT is 
    for VITAL_ACT
    end for;
 end CFG_IOPADN_OUT_VITAL;

 ---- CELL BIBUF_F_2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_2 :  entity is TRUE;
 end BIBUF_F_2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_2_VITAL of BIBUF_F_2 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_2_VITAL;



 ---- CELL BIBUF_F_2D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_2D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_2D :  entity is TRUE;
 end BIBUF_F_2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_2D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_2D_VITAL of BIBUF_F_2D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_2D_VITAL;



 ---- CELL BIBUF_F_2U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_2U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_2U :  entity is TRUE;
 end BIBUF_F_2U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_2U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_2U_VITAL of BIBUF_F_2U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_2U_VITAL;



 ---- CELL BIBUF_F_4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_4 :  entity is TRUE;
 end BIBUF_F_4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_4_VITAL of BIBUF_F_4 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_4_VITAL;



 ---- CELL BIBUF_F_4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_4D :  entity is TRUE;
 end BIBUF_F_4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_4D_VITAL of BIBUF_F_4D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_4D_VITAL;



 ---- CELL BIBUF_F_4U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_4U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_4U :  entity is TRUE;
 end BIBUF_F_4U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_4U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_4U_VITAL of BIBUF_F_4U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_4U_VITAL;



 ---- CELL BIBUF_F_6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_6 :  entity is TRUE;
 end BIBUF_F_6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_6_VITAL of BIBUF_F_6 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_6_VITAL;



 ---- CELL BIBUF_F_6D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_6D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_6D :  entity is TRUE;
 end BIBUF_F_6D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_6D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_6D_VITAL of BIBUF_F_6D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_6D_VITAL;



 ---- CELL BIBUF_F_6U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_F_6U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_F_6U :  entity is TRUE;
 end BIBUF_F_6U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_F_6U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_F_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_F_6U_VITAL of BIBUF_F_6U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_F_6U_VITAL;



 ---- CELL BIBUF_S_2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_2 :  entity is TRUE;
 end BIBUF_S_2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_2_VITAL of BIBUF_S_2 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_2_VITAL;



 ---- CELL BIBUF_S_2D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_2D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_2D :  entity is TRUE;
 end BIBUF_S_2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_2D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_2D_VITAL of BIBUF_S_2D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_2D_VITAL;



 ---- CELL BIBUF_S_2U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_2U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_2U :  entity is TRUE;
 end BIBUF_S_2U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_2U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_2U_VITAL of BIBUF_S_2U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_2U_VITAL;



 ---- CELL BIBUF_S_4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_4 :  entity is TRUE;
 end BIBUF_S_4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_4_VITAL of BIBUF_S_4 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_4_VITAL;



 ---- CELL BIBUF_S_4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_4D :  entity is TRUE;
 end BIBUF_S_4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_4D_VITAL of BIBUF_S_4D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_4D_VITAL;



 ---- CELL BIBUF_S_4U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_4U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_4U :  entity is TRUE;
 end BIBUF_S_4U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_4U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_4U_VITAL of BIBUF_S_4U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_4U_VITAL;



 ---- CELL BIBUF_S_6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_6 :  entity is TRUE;
 end BIBUF_S_6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_6_VITAL of BIBUF_S_6 is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_6_VITAL;



 ---- CELL BIBUF_S_6D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_6D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_6D :  entity is TRUE;
 end BIBUF_S_6D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_6D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_6D_VITAL of BIBUF_S_6D is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_6D_VITAL;



 ---- CELL BIBUF_S_6U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BIBUF_S_6U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BIBUF_S_6U :  entity is TRUE;
 end BIBUF_S_6U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BIBUF_S_6U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/BIBUF_S_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BIBUF_S_6U_VITAL of BIBUF_S_6U is 
    for VITAL_ACT
    end for;
 end CFG_BIBUF_S_6U_VITAL;



 ---- CELL OUTBUF_F_2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_2 :  entity is TRUE;
 end OUTBUF_F_2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_2_VITAL of OUTBUF_F_2 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_2_VITAL;



 ---- CELL OUTBUF_F_4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_4 :  entity is TRUE;
 end OUTBUF_F_4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_4_VITAL of OUTBUF_F_4 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_4_VITAL;



 ---- CELL OUTBUF_F_6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_F_6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_F_6 :  entity is TRUE;
 end OUTBUF_F_6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_F_6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_F_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_F_6_VITAL of OUTBUF_F_6 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_F_6_VITAL;



 ---- CELL OUTBUF_S_2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_2 :  entity is TRUE;
 end OUTBUF_S_2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_2_VITAL of OUTBUF_S_2 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_2_VITAL;



 ---- CELL OUTBUF_S_4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_4 :  entity is TRUE;
 end OUTBUF_S_4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_4_VITAL of OUTBUF_S_4 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_4_VITAL;



 ---- CELL OUTBUF_S_6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OUTBUF_S_6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OUTBUF_S_6 :  entity is TRUE;
 end OUTBUF_S_6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of OUTBUF_S_6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/OUTBUF_S_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(D_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OUTBUF_S_6_VITAL of OUTBUF_S_6 is 
    for VITAL_ACT
    end for;
 end CFG_OUTBUF_S_6_VITAL;



 ---- CELL TRIBUFF_F_2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_2 :  entity is TRUE;
 end TRIBUFF_F_2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_2_VITAL of TRIBUFF_F_2 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_2_VITAL;



 ---- CELL TRIBUFF_F_2D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_2D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_2D :  entity is TRUE;
 end TRIBUFF_F_2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_2D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_2D_VITAL of TRIBUFF_F_2D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_2D_VITAL;



 ---- CELL TRIBUFF_F_2U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_2U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_2U :  entity is TRUE;
 end TRIBUFF_F_2U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_2U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_2U_VITAL of TRIBUFF_F_2U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_2U_VITAL;



 ---- CELL TRIBUFF_F_4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_4 :  entity is TRUE;
 end TRIBUFF_F_4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_4_VITAL of TRIBUFF_F_4 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_4_VITAL;



 ---- CELL TRIBUFF_F_4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_4D :  entity is TRUE;
 end TRIBUFF_F_4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_4D_VITAL of TRIBUFF_F_4D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_4D_VITAL;



 ---- CELL TRIBUFF_F_4U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_4U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_4U :  entity is TRUE;
 end TRIBUFF_F_4U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_4U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_4U_VITAL of TRIBUFF_F_4U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_4U_VITAL;



 ---- CELL TRIBUFF_F_6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_6 :  entity is TRUE;
 end TRIBUFF_F_6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_6_VITAL of TRIBUFF_F_6 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_6_VITAL;



 ---- CELL TRIBUFF_F_6D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_6D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_6D :  entity is TRUE;
 end TRIBUFF_F_6D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_6D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_6D_VITAL of TRIBUFF_F_6D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_6D_VITAL;



 ---- CELL TRIBUFF_F_6U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_F_6U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_F_6U :  entity is TRUE;
 end TRIBUFF_F_6U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_F_6U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_F_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_F_6U_VITAL of TRIBUFF_F_6U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_F_6U_VITAL;



 ---- CELL TRIBUFF_S_2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_2 :  entity is TRUE;
 end TRIBUFF_S_2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

        begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_2",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_2_VITAL of TRIBUFF_S_2 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_2_VITAL;



 ---- CELL TRIBUFF_S_2D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_2D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_2D :  entity is TRUE;
 end TRIBUFF_S_2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_2D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_2D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_2D_VITAL of TRIBUFF_S_2D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_2D_VITAL;



 ---- CELL TRIBUFF_S_2U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_2U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_2U :  entity is TRUE;
 end TRIBUFF_S_2U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_2U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_2U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_2U_VITAL of TRIBUFF_S_2U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_2U_VITAL;



 ---- CELL TRIBUFF_S_4 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_4 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_4 :  entity is TRUE;
 end TRIBUFF_S_4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_4 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_4",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_4_VITAL of TRIBUFF_S_4 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_4_VITAL;



 ---- CELL TRIBUFF_S_4D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_4D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_4D :  entity is TRUE;
 end TRIBUFF_S_4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_4D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_4D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_4D_VITAL of TRIBUFF_S_4D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_4D_VITAL;



 ---- CELL TRIBUFF_S_4U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_4U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_4U :  entity is TRUE;
 end TRIBUFF_S_4U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_4U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_4U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_4U_VITAL of TRIBUFF_S_4U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_4U_VITAL;



 ---- CELL TRIBUFF_S_6 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_6 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_6 :  entity is TRUE;
 end TRIBUFF_S_6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_6 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_6",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_6_VITAL of TRIBUFF_S_6 is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_6_VITAL;



 ---- CELL TRIBUFF_S_6D ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_6D is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_6D :  entity is TRUE;
 end TRIBUFF_S_6D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_6D is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_6D",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01LWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_6D_VITAL of TRIBUFF_S_6D is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_6D_VITAL;



 ---- CELL TRIBUFF_S_6U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity TRIBUFF_S_6U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of TRIBUFF_S_6U :  entity is TRUE;
 end TRIBUFF_S_6U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of TRIBUFF_S_6U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/TRIBUFF_S_6U",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_TRIBUFF_S_6U_VITAL of TRIBUFF_S_6U is 
    for VITAL_ACT
    end for;
 end CFG_TRIBUFF_S_6U_VITAL;



 ---- CELL BUFD ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BUFD is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BUFD :  entity is TRUE;
 end BUFD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of BUFD is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BUFD_VITAL of BUFD is 
    for VITAL_ACT
    end for;
 end CFG_BUFD_VITAL;



 ---- CELL INVD ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INVD is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INVD :  entity is TRUE;
 end INVD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of INVD is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INVD_VITAL of INVD is 
    for VITAL_ACT
    end for;
 end CFG_INVD_VITAL;



 ---- CELL IOIN_IR ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IR is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_IR :  entity is TRUE;
 end IOIN_IR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IR is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	  VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, ICLK_ipd)

	-- timing check results
	VARIABLE Tviol_YIN_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_YIN_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_ICLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_ICLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE ICLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE YIN_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_YIN_ICLK_posedge,
	 TimingData		=> Tmkr_YIN_ICLK_posedge,
	 TestSignal		=> YIN_ipd,
	 TestSignalName		=> "YIN",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName	        => "ICLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_YIN_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_YIN_ICLK_negedge_posedge,
	 HoldHigh		=> thold_YIN_ICLK_posedge_posedge,
	 HoldLow		=> thold_YIN_ICLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOIN_IR",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_ICLK,
	 PeriodData		=> PInfo_ICLK,
	 TestSignal		=> ICLK_ipd,
	 TestSignalName		=> "ICLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_ICLK_posedge,
	 PulseWidthLow		=> tpw_ICLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "IOIN_IR",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_YIN_ICLK_posedge or 
	 Pviol_ICLK;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Y,
	 GlitchData => Y_GlitchData,
	 OutSignalName => "Y",
	 OutTemp => Y_zd,
	 Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOIN_IR_VITAL of IOIN_IR is
   for VITAL_ACT
   end for;
end CFG_IOIN_IR_VITAL;



 ---- CELL IOIN_IRE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_IRE is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_ICLK_Y		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_ICE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		ICE		:   in    STD_ULOGIC;
		ICLK		:   in    STD_ULOGIC;
		YIN		:  in    STD_ULOGIC;
		Y		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_IRE :  entity is TRUE;
 end IOIN_IRE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_IRE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICE_ipd  : STD_ULOGIC := 'X';
	SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
	  VitalWireDelay (ICE_ipd,ICE, tipd_ICE);
	  VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, ICE_ipd,ICLK_ipd)

	-- timing check results
	VARIABLE Tviol_YIN_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_YIN_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_ICE_ICLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_ICE_ICLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_ICLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_ICLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE ICE_delayed	: STD_ULOGIC := 'X';
	VARIABLE ICLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE YIN_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_YIN_ICLK_posedge,
	 TimingData		=> Tmkr_YIN_ICLK_posedge,
	 TestSignal		=> YIN_ipd,
	 TestSignalName		=> "YIN",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName	        => "ICLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_YIN_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_YIN_ICLK_negedge_posedge,
	 HoldHigh		=> thold_YIN_ICLK_posedge_posedge,
	 HoldLow		=> thold_YIN_ICLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((ICE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOIN_IRE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_ICE_ICLK_posedge,
	 TimingData		=> Tmkr_ICE_ICLK_posedge,
	 TestSignal		=> ICE_ipd,
	 TestSignalName		=> "ICE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> ICLK_ipd,
	 RefSignalName		=> "ICLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_ICE_ICLK_posedge_posedge,
	 SetupLow		=> tsetup_ICE_ICLK_negedge_posedge,
	 HoldHigh		=> thold_ICE_ICLK_posedge_posedge,
	 HoldLow		=> thold_ICE_ICLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOIN_IRE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_ICLK,
	 PeriodData		=> PInfo_ICLK,
	 TestSignal		=> ICLK_ipd,
	 TestSignalName		=> "ICLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_ICLK_posedge,
	 PulseWidthLow		=> tpw_ICLK_negedge,
	 CheckEnabled		=> TRUE,
	 HeaderMsg		=> InstancePath & "IOIN_IRE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_YIN_ICLK_posedge or 
	 Tviol_ICE_ICLK_posedge or 
	 Pviol_ICLK;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Y,
	 GlitchData => Y_GlitchData,
	 OutSignalName => "Y",
	 OutTemp => Y_zd,
	 Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOIN_IRE_VITAL of IOIN_IRE is
   for VITAL_ACT
   end for;
end CFG_IOIN_IRE_VITAL;



 ---- CELL IOTRI_OB_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_ER is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OB_ER :  entity is TRUE;
 end IOTRI_OB_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_ER is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_E_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS EOUT_zd : STD_LOGIC is Results(1);
	ALIAS DOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_OCLK_posedge,
	 TimingData		=> Tmkr_E_OCLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_E_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_E_OCLK_negedge_posedge,
	 HoldHigh		=> thold_E_OCLK_posedge_posedge,
	 HoldLow		=> thold_E_OCLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OB_ER",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ER",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_E_OCLK_posedge or 
	 Pviol_OCLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
    --- combinatorial output logic. 
   DOUT_zd :=  D_ipd ;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (
	         0 => (D_ipd'last_event, tpd_D_DOUT, true),
	           1 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OB_ER_VITAL of IOTRI_OB_ER is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OB_ER_VITAL;



 ---- CELL IOTRI_OB_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OB_ERE is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_DOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OB_ERE :  entity is TRUE;
 end IOTRI_OB_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OB_ERE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (OCE_ipd,OCE, tipd_OCE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_E_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_E_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_OCE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_OCE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCE_delayed	: STD_ULOGIC := 'X';
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE E_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS EOUT_zd : STD_LOGIC is Results(1);
	ALIAS DOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_E_OCLK_posedge,
	 TimingData		=> Tmkr_E_OCLK_posedge,
	 TestSignal		=> E_ipd,
	 TestSignalName		=> "E",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_E_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_E_OCLK_negedge_posedge,
	 HoldHigh		=> thold_E_OCLK_posedge_posedge,
	 HoldLow		=> thold_E_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((OCE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OB_ERE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_OCE_OCLK_posedge,
	 TimingData		=> Tmkr_OCE_OCLK_posedge,
	 TestSignal		=> OCE_ipd,
	 TestSignalName		=> "OCE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_OCE_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_OCE_OCLK_negedge_posedge,
	 HoldHigh		=> thold_OCE_OCLK_posedge_posedge,
	 HoldLow		=> thold_OCE_OCLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_OB_ERE",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_E_OCLK_posedge or 
	 Tviol_OCE_OCLK_posedge or 
	 Pviol_OCLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
    --- combinatorial output logic. 
   DOUT_zd :=  D_ipd ;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (
	         0 => (D_ipd'last_event, tpd_D_DOUT, true),
	           1 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OB_ERE_VITAL of IOTRI_OB_ERE is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OB_ERE_VITAL;



 ---- CELL IOTRI_OR_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OR_EB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OR_EB :  entity is TRUE;
 end IOTRI_OR_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OR_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_OCLK_posedge,
	 TimingData		=> Tmkr_D_OCLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_D_OCLK_negedge_posedge,
	 HoldHigh		=> thold_D_OCLK_posedge_posedge,
	 HoldLow		=> thold_D_OCLK_negedge_posedge,
	 CheckEnabled		=>  TRUE, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_OR_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_OR_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_OCLK_posedge or 
	 Pviol_OCLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
    --- combinatorial output logic. 
   EOUT_zd :=  E_ipd ;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (
	         0 => (E_ipd'last_event, tpd_E_EOUT, true),
	           1 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OR_EB_VITAL of IOTRI_OR_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OR_EB_VITAL;



 ---- CELL IOTRI_ORE_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_ORE_EB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_DOUT		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT		:   VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_OCE		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		OCE		:   in    STD_ULOGIC;
		OCLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		E		:  in    STD_ULOGIC;
		DOUT		:  out    STD_ULOGIC;
		EOUT		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_ORE_EB :  entity is TRUE;
 end IOTRI_ORE_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_ORE_EB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
	SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (E_ipd, E, tipd_E);
	  VitalWireDelay (OCE_ipd,OCE, tipd_OCE);
	  VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCE_ipd,OCLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_OCE_OCLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_OCE_OCLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_OCLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_OCLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE OCE_delayed	: STD_ULOGIC := 'X';
	VARIABLE OCLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS DOUT_zd : STD_LOGIC is Results(1);
	ALIAS EOUT_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
	VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_OCLK_posedge,
	 TimingData		=> Tmkr_D_OCLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName	        => "OCLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_D_OCLK_negedge_posedge,
	 HoldHigh		=> thold_D_OCLK_posedge_posedge,
	 HoldLow		=> thold_D_OCLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((OCE_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/IOTRI_ORE_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalSetupHoldCheck (
	 Violation		=> Tviol_OCE_OCLK_posedge,
	 TimingData		=> Tmkr_OCE_OCLK_posedge,
	 TestSignal		=> OCE_ipd,
	 TestSignalName		=> "OCE",
	 TestDelay		=> 0 ns,
	 RefSignal		=> OCLK_ipd,
	 RefSignalName		=> "OCLK",
	 RefDelay 		=> 0 ns,
	 SetupHigh		=> tsetup_OCE_OCLK_posedge_posedge,
	 SetupLow		=> tsetup_OCE_OCLK_negedge_posedge,
	 HoldHigh		=> thold_OCE_OCLK_posedge_posedge,
	 HoldLow		=> thold_OCE_OCLK_negedge_posedge,
	 CheckEnabled		=>  TRUE,	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "IOTRI_ORE_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_OCLK,
	 PeriodData		=> PInfo_OCLK,
	 TestSignal		=> OCLK_ipd,
	 TestSignalName		=> "OCLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_OCLK_posedge,
	 PulseWidthLow		=> tpw_OCLK_negedge,
	 CheckEnabled		=>TRUE,
	 HeaderMsg		=> InstancePath & "IOTRI_ORE_EB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_OCLK_posedge or 
	 Tviol_OCE_OCLK_posedge or 
	 Pviol_OCLK;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
    --- combinatorial output logic. 
   EOUT_zd :=  E_ipd ;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => DOUT,
	 GlitchData => DOUT_GlitchData,
	 OutSignalName => "DOUT",
	 OutTemp => DOUT_zd,
	 Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

	VitalPathDelay01 (
	 OutSignal => EOUT,
	 GlitchData => EOUT_GlitchData,
	 OutSignalName => "EOUT",
	 OutTemp => EOUT_zd,
	 Paths => (
	         0 => (E_ipd'last_event, tpd_E_EOUT, true),
	           1 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_ORE_EB_VITAL of IOTRI_ORE_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_ORE_EB_VITAL;



 ---- CELL IOTRI_ORE_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_ORE_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_ORE_ERE :  entity is TRUE;
 end IOTRI_ORE_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_ORE_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, OCLK_ipd, OCE_ipd, D_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_ORE_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_D_OCLK_posedge ;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOTRI_ORE_ERE_VITAL of IOTRI_ORE_ERE is
   for VITAL_ACT
   end for;
end CFG_IOTRI_ORE_ERE_VITAL;



 ---- CELL IOTRI_OR_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OR_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOTRI_OR_ER :  entity is TRUE;
 end IOTRI_OR_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OR_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, OCLK_ipd, D_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOTRI_OR_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOTRI_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_D_OCLK_posedge ;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OR_ER_VITAL of IOTRI_OR_ER is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OR_ER_VITAL;



 ---- CELL IOBI_IB_OB_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_ER :  entity is TRUE;
 end IOBI_IB_OB_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, YIN_ipd, E_ipd, OCLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);
   ALIAS EOUT_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK;

        DOUT_zd :=TO_X01(D_ipd);

        Y_zd :=TO_X01(YIN_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OB_ER_VITAL of IOBI_IB_OB_ER is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OB_ER_VITAL;



 ---- CELL IOBI_IB_OB_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OB_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OB_ERE :  entity is TRUE;
 end IOBI_IB_OB_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OB_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, YIN_ipd, E_ipd, OCLK_ipd, OCE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);
   ALIAS EOUT_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OB_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

        Y_zd :=TO_X01(YIN_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;



   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OB_ERE_VITAL of IOBI_IB_OB_ERE is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OB_ERE_VITAL;



 ---- CELL IOBI_IB_OR_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OR_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_Yin_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_Yin :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                Yin         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OR_EB :  entity is TRUE;
 end IOBI_IB_OR_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OR_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL Yin_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (Yin_ipd, Yin, tipd_Yin);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, Yin_ipd, D_ipd, OCLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Yin_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);
   ALIAS DOUT_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OR_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OR_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK;

        EOUT_zd :=TO_X01(E_ipd);

        Y_zd :=TO_X01(Yin_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (Yin_ipd'last_event, tpd_Yin_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OR_EB_VITAL of IOBI_IB_OR_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OR_EB_VITAL;



 ---- CELL IOBI_IB_ORE_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_ORE_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_ORE_EB :  entity is TRUE;
 end IOBI_IB_ORE_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_ORE_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, YIN_ipd, D_ipd, OCLK_ipd, OCE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);
   ALIAS DOUT_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORE_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

        Y_zd :=TO_X01(YIN_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_ORE_EB_VITAL of IOBI_IB_ORE_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_ORE_EB_VITAL;



 ---- CELL IOBI_IB_OR_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_OR_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                YIN         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_OR_ER :  entity is TRUE;
 end IOBI_IB_OR_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_OR_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, D_ipd, OCLK_ipd, E_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS EOUT_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE Y_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_OR_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_E_OCLK_posedge ;

        Y_zd :=TO_X01(YIN_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_OR_ER_VITAL of IOBI_IB_OR_ER is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_OR_ER_VITAL;



 ---- CELL IOBI_IB_ORE_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IB_ORE_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_YIN_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                YIN         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                Y                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IB_ORE_ERE :  entity is TRUE;
 end IOBI_IB_ORE_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IB_ORE_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, D_ipd, OCLK_ipd, OCE_ipd, E_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS EOUT_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE Y_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IB_ORE_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IB_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_E_OCLK_posedge ;

        Y_zd :=TO_X01(YIN_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (YIN_ipd'last_event, tpd_YIN_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IB_ORE_ERE_VITAL of IOBI_IB_ORE_ERE is
   for VITAL_ACT
   end for;
end CFG_IOBI_IB_ORE_ERE_VITAL;



 ---- CELL IOBI_IR_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_OB_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_OB_EB :  entity is TRUE;
 end IOBI_IR_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_OB_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        DOUT_zd :=TO_X01(D_ipd);

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_OB_EB_VITAL of IOBI_IR_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_OB_EB_VITAL;



 ---- CELL IOBI_IRE_OB_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_OB_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_OB_EB :  entity is TRUE;
 end IOBI_IRE_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_OB_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OB_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_OB_EB_VITAL of IOBI_IRE_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_OB_EB_VITAL;



 ---- CELL IOBI_IR_OB_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_OB_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_OB_ER :  entity is TRUE;
 end IOBI_IR_OB_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_OB_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OB_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OB_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OB_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OB_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_OB_ER_VITAL of IOBI_IR_OB_ER is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_OB_ER_VITAL;



 ---- CELL IOBI_IRE_OB_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_OB_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_OB_ER :  entity is TRUE;
 end IOBI_IRE_OB_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_OB_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OB_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OB_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_OB_ER_VITAL of IOBI_IRE_OB_ER is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_OB_ER_VITAL;



 ---- CELL IOBI_IR_OB_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_OB_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_OB_ERE :  entity is TRUE;
 end IOBI_IR_OB_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_OB_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, OCE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OB_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OB_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_OB_ERE_VITAL of IOBI_IR_OB_ERE is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_OB_ERE_VITAL;



 ---- CELL IOBI_IRE_OB_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_OB_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_D_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                D         : in    STD_ULOGIC;
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_OB_ERE :  entity is TRUE;
 end IOBI_IRE_OB_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_OB_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, OCLK_ipd, OCE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS DOUT_zd : STD_LOGIC is Results(1);
   ALIAS EOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OB_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OB_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OB_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        DOUT_zd :=TO_X01(D_ipd);

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_OB_ERE_VITAL of IOBI_IRE_OB_ERE is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_OB_ERE_VITAL;



 ---- CELL IOBI_IR_OR_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_OR_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_OR_EB :  entity is TRUE;
 end IOBI_IR_OR_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_OR_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);

   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OR_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OR_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OR_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OR_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_OR_EB_VITAL of IOBI_IR_OR_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_OR_EB_VITAL;



 ---- CELL IOBI_IRE_OR_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_OR_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_OR_EB :  entity is TRUE;
 end IOBI_IRE_OR_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_OR_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OR_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OR_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_OR_EB_VITAL of IOBI_IRE_OR_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_OR_EB_VITAL;



 ---- CELL IOBI_IR_ORE_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_ORE_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_ORE_EB :  entity is TRUE;
 end IOBI_IR_ORE_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_ORE_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, OCE_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_ORE_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_ORE_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_ORE_EB_VITAL of IOBI_IR_ORE_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_ORE_EB_VITAL;



 ---- CELL IOBI_IRE_ORE_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_ORE_EB is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_E_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_ORE_EB :  entity is TRUE;
 end IOBI_IRE_ORE_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_ORE_EB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, D_ipd, OCLK_ipd, OCE_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);

   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_ORE_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_ORE_EB",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_EB",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_D_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

        EOUT_zd :=TO_X01(E_ipd);

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_ORE_EB_VITAL of IOBI_IRE_ORE_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_ORE_EB_VITAL;



 ---- CELL IOBI_IR_OR_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_OR_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_OR_ER :  entity is TRUE;
 end IOBI_IR_OR_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_OR_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, OCLK_ipd, D_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_3  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OR_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_OR_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_D_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_3,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_OR_ER_VITAL of IOBI_IR_OR_ER is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_OR_ER_VITAL;



 ---- CELL IOBI_IR_ORE_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IR_ORE_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IR_ORE_ERE :  entity is TRUE;
 end IOBI_IR_ORE_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IR_ORE_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, OCLK_ipd, OCE_ipd, D_ipd, YIN_ipd, ICLK_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_3  : STD_LOGIC_VECTOR(0 to 6);

   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_ORE_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IR_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IR_ORE_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_D_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_3,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed, '0', '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IR_ORE_ERE_VITAL of IOBI_IR_ORE_ERE is
   for VITAL_ACT
   end for;
end CFG_IOBI_IR_ORE_ERE_VITAL;



 ---- CELL IOBI_IRE_OR_ER ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_OR_ER is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_OR_ER :  entity is TRUE;
 end IOBI_IRE_OR_ER;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_OR_ER is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, OCLK_ipd, D_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_3  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OR_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_OR_ER",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_OR_ER",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_D_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed, '0', '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed, '0', '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_3,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_OR_ER_VITAL of IOBI_IRE_OR_ER is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_OR_ER_VITAL;



 ---- CELL IOBI_IRE_ORE_ERE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_IRE_ORE_ERE is
	generic(
		TimingChecksOn: Boolean := True;
		InstancePath: STRING := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_OCLK_EOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_OCLK_DOUT	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_ICLK_Y	:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_E_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_E_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_OCLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_OCLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_OCE_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_OCE_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_D_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_D_OCLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_D_OCLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_YIN_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tpw_ICLK_posedge	:  VitalDelayType := 0.000 ns;
		tpw_ICLK_negedge	:  VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
		tsetup_ICE_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_posedge_posedge	:   VitalDelayType := 0.000 ns;
		thold_ICE_ICLK_negedge_posedge       :   VitalDelayType := 0.000 ns;
		tipd_E :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_OCE :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_YIN :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICLK :   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_ICE :   VitalDelayType01 := (0.000 ns, 0.000 ns));
    port(
                E         : in    STD_ULOGIC;
                OCLK         : in    STD_ULOGIC;
                OCE         : in    STD_ULOGIC;
                D         : in    STD_ULOGIC;
                YIN         : in    STD_ULOGIC;
                ICLK         : in    STD_ULOGIC;
                ICE         : in    STD_ULOGIC;
                EOUT                : out    STD_ULOGIC;
                DOUT                : out    STD_ULOGIC;
                Y                : out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBI_IRE_ORE_ERE :  entity is TRUE;
 end IOBI_IRE_ORE_ERE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_IRE_ORE_ERE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL E_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL OCE_ipd  : STD_ULOGIC := 'X';
   SIGNAL D_ipd  : STD_ULOGIC := 'X';
   SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICLK_ipd  : STD_ULOGIC := 'X';
   SIGNAL ICE_ipd  : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (OCLK_ipd, OCLK, tipd_OCLK);
   VitalWireDelay (OCE_ipd, OCE, tipd_OCE);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
   VitalWireDelay (ICLK_ipd, ICLK, tipd_ICLK);
   VitalWireDelay (ICE_ipd, ICE, tipd_ICE);
   end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (E_ipd, OCLK_ipd, OCE_ipd, D_ipd, YIN_ipd, ICLK_ipd, ICE_ipd)


   VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_E_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_OCLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_OCLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_OCE_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_OCE_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_OCLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_D_OCLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_YIN_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_ICLK    : STD_ULOGIC := '0';
   VARIABLE PInfo_ICLK    : VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Tviol_ICE_ICLK_posedge         : STD_ULOGIC := '0';
   VARIABLE Tmkr_ICE_ICLK_posedge         : VitalTimingDataType := VitalTimingDataInit;

   -- functionality results
   VARIABLE Violation      : STD_ULOGIC := '0';
   VARIABLE PrevData_Q_1  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_2  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE PrevData_Q_3  : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE E_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE OCE_delayed       : STD_ULOGIC := 'X';
   VARIABLE D_delayed       : STD_ULOGIC := 'X';
   VARIABLE YIN_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICLK_delayed       : STD_ULOGIC := 'X';
   VARIABLE ICE_delayed       : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3)  := (others => 'X');
   ALIAS EOUT_zd : STD_LOGIC is Results(1);
   ALIAS DOUT_zd : STD_LOGIC is Results(2);
   ALIAS Y_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE EOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
   VARIABLE Y_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
  VitalSetupHoldCheck (
   Violation              => Tviol_E_OCLK_posedge,
   TimingData             => Tmkr_E_OCLK_posedge,
   TestSignal             => E_ipd,
   TestSignalName         => "E",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_E_OCLK_posedge_posedge,
   SetupLow               => tsetup_E_OCLK_negedge_posedge,
   HoldHigh              => thold_E_OCLK_posedge_posedge,
   HoldLow                => thold_E_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_OCLK,
    PeriodData             => PInfo_OCLK,
    TestSignal             => OCLK_ipd,
    TestSignalName         => "OCLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_OCLK_posedge,
    PulseWidthLow          => tpw_OCLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_ORE_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_OCE_OCLK_posedge,
   TimingData             => Tmkr_OCE_OCLK_posedge,
   TestSignal             => OCE_ipd,
   TestSignalName         => "OCE",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_OCE_OCLK_posedge_posedge,
   SetupLow               => tsetup_OCE_OCLK_negedge_posedge,
   HoldHigh              => thold_OCE_OCLK_posedge_posedge,
   HoldLow                => thold_OCE_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_D_OCLK_posedge,
   TimingData             => Tmkr_D_OCLK_posedge,
   TestSignal             => D_ipd,
   TestSignalName         => "D",
   TestDelay              => 0 ns,
   RefSignal              => OCLK_ipd,
   RefSignalName          => "OCLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_D_OCLK_posedge_posedge,
   SetupLow               => tsetup_D_OCLK_negedge_posedge,
   HoldHigh              => thold_D_OCLK_posedge_posedge,
   HoldLow                => thold_D_OCLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_YIN_ICLK_posedge,
   TimingData             => Tmkr_YIN_ICLK_posedge,
   TestSignal             => YIN_ipd,
   TestSignalName         => "YIN",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
   SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
   HoldHigh              => thold_YIN_ICLK_posedge_posedge,
   HoldLow                => thold_YIN_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   VitalPeriodPulseCheck (
    Violation              => Pviol_ICLK,
    PeriodData             => PInfo_ICLK,
    TestSignal             => ICLK_ipd,
    TestSignalName         => "ICLK",
    TestDelay              => 0 ns,
    Period         => 0 ns,
    PulseWidthHigh => tpw_ICLK_posedge,
    PulseWidthLow          => tpw_ICLK_negedge,
    CheckEnabled           => TRUE,
    HeaderMsg              => InstancePath & "IOBI_IRE_ORE_ERE",
    Xon            => Xon,
    MsgOn          => MsgOn,
    MsgSeverity            => WARNING);

  VitalSetupHoldCheck (
   Violation              => Tviol_ICE_ICLK_posedge,
   TimingData             => Tmkr_ICE_ICLK_posedge,
   TestSignal             => ICE_ipd,
   TestSignalName         => "ICE",
   TestDelay              => 0 ns,
   RefSignal              => ICLK_ipd,
   RefSignalName          => "ICLK",
   RefDelay               => 0 ns,
   SetupHigh              => tsetup_ICE_ICLK_posedge_posedge,
   SetupLow               => tsetup_ICE_ICLK_negedge_posedge,
   HoldHigh              => thold_ICE_ICLK_posedge_posedge,
   HoldLow                => thold_ICE_ICLK_negedge_posedge,
   CheckEnabled           => TRUE,
   RefTransition          => 'R',
   HeaderMsg              => InstancePath & "/IOBI_IRE_ORE_ERE",
   Xon            => Xon,
   MsgOn          => MsgOn,
   MsgSeverity    => WARNING);

   end if;

   -------------------------
   --  Functionality Section
   -------------------------

   Violation :=  Tviol_E_OCLK_posedge  or Pviol_OCLK or Tviol_OCE_OCLK_posedge  or Tviol_D_OCLK_posedge  or Tviol_YIN_ICLK_posedge  or Pviol_ICLK or Tviol_ICE_ICLK_posedge ;

  VitalStateTable(
   Result => EOUT_zd,
   PreviousDataIn => PrevData_Q_1,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, EOUT_zd, E_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   EOUT_zd := Violation XOR EOUT_zd;
   E_delayed := E_ipd;

  VitalStateTable(
   Result => DOUT_zd,
   PreviousDataIn => PrevData_Q_2,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', OCLK_delayed, DOUT_zd, D_delayed,  (NOT OCE_delayed), '1', OCLK_ipd));
   DOUT_zd := Violation XOR DOUT_zd;
   D_delayed := D_ipd;
   OCE_delayed := OCE_ipd;
   OCLK_delayed := OCLK_ipd;

  VitalStateTable(
   Result => Y_zd,
   PreviousDataIn => PrevData_Q_3,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', ICLK_delayed, Y_zd, YIN_delayed,  (NOT ICE_delayed), '1', ICLK_ipd));
   Y_zd := Violation XOR Y_zd;
   YIN_delayed := YIN_ipd;
   ICE_delayed := ICE_ipd;
   ICLK_delayed := ICLK_ipd;


   ----------------------
   --  Path Delay Section
   ----------------------
   VitalPathDelay01 (
    OutSignal => EOUT,
    GlitchData => EOUT_GlitchData,
    OutSignalName => "EOUT",
    OutTemp => EOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => DOUT,
    GlitchData => DOUT_GlitchData,
    OutSignalName => "DOUT",
    OutTemp => DOUT_zd,
    Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);

   VitalPathDelay01 (
    OutSignal => Y,
    GlitchData => Y_GlitchData,
    OutSignalName => "Y",
    OutTemp => Y_zd,
    Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_Y, true)),
    Mode => OnDetect,
    Xon => Xon,
    MsgOn => MsgOn,
    MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_IOBI_IRE_ORE_ERE_VITAL of IOBI_IRE_ORE_ERE is
   for VITAL_ACT
   end for;
end CFG_IOBI_IRE_ORE_ERE_VITAL;



 ---- CELL CLKIO ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKIO is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKIO :  entity is TRUE;
 end CLKIO;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKIO is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKIO_VITAL of CLKIO is 
    for VITAL_ACT
    end for;
 end CFG_CLKIO_VITAL;


 ---- CELL CLKBIBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity CLKBIBUF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: STRING :="*";
		MsgOn: Boolean := True;

                tpw_D_posedge           : VitalDelayType := 0.000 ns;
                tpw_D_negedge           : VitalDelayType := 0.000 ns;
                tpw_E_posedge           : VitalDelayType := 0.000 ns;
                tpw_E_negedge           : VitalDelayType := 0.000 ns;
                tpw_PAD_negedge         : VitalDelayType := 0.000 ns;
                tpw_PAD_posedge         : VitalDelayType := 0.000 ns;

		tpd_D_PAD		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_E_PAD : VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_D_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
			tpd_E_Y			: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_D		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_E		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		D		: in    STD_ULOGIC;
		E		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of CLKBIBUF :  entity is TRUE;
 end CLKBIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of CLKBIBUF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL E_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (E_ipd, E, tipd_E);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)

        -- timing check results
        VARIABLE Pviol_D        : STD_ULOGIC := '0';
        VARIABLE PeriodData_D   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_E        : STD_ULOGIC := '0';
        VARIABLE PeriodData_E   : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_PAD      : STD_ULOGIC := '0';
        VARIABLE PeriodData_PAD : VitalPeriodDataType := VitalPeriodDataInit;



	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

        -- timing check results
        if( TimingChecksOn ) then

            VitalPeriodPulseCheck (
              Violation      => Pviol_PAD,
              PeriodData     => PeriodData_PAD,
              TestSignal     => PAD_ipd,
              TestSignalName => "PAD",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_PAD_posedge,
              PulseWidthLow  => tpw_PAD_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBIBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_D,
              PeriodData     => PeriodData_D,
              TestSignal     => D_ipd,
              TestSignalName => "D",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_D_posedge,
              PulseWidthLow  => tpw_D_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBIBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );


            VitalPeriodPulseCheck (
              Violation      => Pviol_E,
              PeriodData     => PeriodData_E,
              TestSignal     => E_ipd,
              TestSignalName => "E",
              TestDelay      => 0 ns,
              Period         => 0 ns,
              PulseWidthHigh => tpw_E_posedge,
              PulseWidthLow  => tpw_E_negedge,
              CheckEnabled   => TRUE,
              HeaderMsg      => InstancePath &"/CLKBIBUF",
              Xon            => Xon,
              MsgOn          => MsgOn,
              MsgSeverity    => WARNING
            );

        end if;


	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => D_ipd,
                   enable =>(NOT E_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (D_ipd'last_event,VitalExtendToFillDelay(tpd_D_PAD),true),
	             1 => (E_ipd'last_event, tpd_E_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (D_ipd'last_event,tpd_D_Y, true),
	             1 => (E_ipd'last_event,tpd_E_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_CLKBIBUF_VITAL of CLKBIBUF is 
    for VITAL_ACT
    end for;
 end CFG_CLKBIBUF_VITAL;


---- CELL DDR_OUT ----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
 entity DDR_OUT is
  generic (
           TimingChecksOn : Boolean := True;
           InstancePath   : STRING  := "*";
           Xon            : Boolean := False;
           MsgOn          : Boolean := True;

           tpd_CLR_Q                         : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
           tpd_CLK_Q                         : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
           tsetup_DR_CLK_posedge_posedge     : VitalDelayType   := 0.000 ns;
           thold_DR_CLK_posedge_posedge      : VitalDelayType   := 0.000 ns;
           tsetup_DR_CLK_negedge_posedge     : VitalDelayType   := 0.000 ns;
           thold_DR_CLK_negedge_posedge      : VitalDelayType   := 0.000 ns;

           tsetup_DF_CLK_posedge_posedge     : VitalDelayType   := 0.000 ns;
           thold_DF_CLK_posedge_posedge      : VitalDelayType   := 0.000 ns;
           tsetup_DF_CLK_negedge_posedge     : VitalDelayType   := 0.000 ns;
           thold_DF_CLK_negedge_posedge      : VitalDelayType   := 0.000 ns;

           thold_CLR_CLK_negedge_posedge     : VitalDelayType   := 0.000 ns;
           trecovery_CLR_CLK_negedge_posedge : VitalDelayType   := 0.000 ns;
           tperiod_CLK_posedge               : VitalDelayType   := 0.000 ns;
           tpw_CLK_posedge                   : VitalDelayType   := 0.000 ns;
           tpw_CLK_negedge                   : VitalDelayType   := 0.000 ns;
           tpw_CLR_posedge                   : VitalDelayType   := 0.000 ns;
           tipd_DR                           : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
           tipd_DF                           : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
           tipd_CLR                          : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
           tipd_CLK                          : VitalDelayType01 := ( 0.000 ns, 0.000 ns )
          );

  port    (
           CLR : in  STD_ULOGIC;
           CLK : in  STD_ULOGIC;
           DR  : in  STD_ULOGIC;
           DF  : in  STD_ULOGIC;
           Q   : out STD_ULOGIC
          );

  attribute VITAL_LEVEL0 of DDR_OUT :  entity is TRUE;
end DDR_OUT;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DDR_OUT is
  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

  SIGNAL DR_ipd  : STD_ULOGIC := 'X';
  SIGNAL DF_ipd  : STD_ULOGIC := 'X';
  SIGNAL CLR_ipd : STD_ULOGIC := 'X';
  SIGNAL CLK_ipd : STD_ULOGIC := 'X';

  begin

    ---------------------
    --  INPUT PATH DELAYs
    ---------------------
    WireDelay : block
      begin
        VitalWireDelay ( DR_ipd,  DR,  tipd_DR );
        VitalWireDelay ( DF_ipd,  DF,  tipd_DF );
        VitalWireDelay ( CLR_ipd, CLR, tipd_CLR );
        VitalWireDelay ( CLK_ipd, CLK, tipd_CLK );
    end block;

    --------------------
    --  BEHAVIOR SECTION
    --------------------
    VITALBehavior : process ( DR_ipd, DF_ipd, CLR_ipd, CLK_ipd )

      -- timing check results
      VARIABLE Tviol_DR_CLK_posedge  : STD_ULOGIC := '0';
      VARIABLE Tmkr_DR_CLK_posedge   : VitalTimingDataType := VitalTimingDataInit;
      VARIABLE Tviol_DF_CLK_posedge  : STD_ULOGIC := '0';
      VARIABLE Tmkr_DF_CLK_posedge   : VitalTimingDataType := VitalTimingDataInit;

      VARIABLE Tviol_CLR_CLK_posedge : STD_ULOGIC := '0';
      VARIABLE Tmkr_CLR_CLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
      VARIABLE Pviol_CLK             : STD_ULOGIC := '0';
      VARIABLE PInfo_CLK             : VitalPeriodDataType := VitalPeriodDataInit;
      VARIABLE Pviol_CLR             : STD_ULOGIC := '0';
      VARIABLE PInfo_CLR             : VitalPeriodDataType := VitalPeriodDataInit;

      -- functionality results
      VARIABLE Violation    : STD_ULOGIC := '0';
      VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 2);
      VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 2);
      VARIABLE QR_tmp       : STD_ULOGIC := 'X';
      VARIABLE QF_tmp       : STD_ULOGIC := 'X';

      VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');

      ALIAS Q_zd : STD_LOGIC is Results(1);

      -- output glitch detection variables
      VARIABLE Q_GlitchData  : VitalGlitchDataType;

      begin


        ------------------------
        --  Timing Check Section
        ------------------------

        if ( TimingChecksOn ) then
          VitalSetupHoldCheck (
            Violation      => Tviol_DR_CLK_posedge,
            TimingData     => Tmkr_DR_CLK_posedge,
            TestSignal     => DR_ipd,
            TestSignalName => "DR",
            TestDelay      => 0 ns,
            RefSignal      => CLK_ipd,
            RefSignalName  => "CLK",
            RefDelay       => 0 ns,
            SetupHigh      => tsetup_DR_CLK_posedge_posedge,
            SetupLow       => tsetup_DR_CLK_negedge_posedge,
            HoldHigh       => thold_DR_CLK_posedge_posedge,
            HoldLow        => thold_DR_CLK_negedge_posedge,
            CheckEnabled   => TO_X01 (( NOT CLR_ipd )) /= '0',
            RefTransition  => 'R',
            HeaderMsg      => InstancePath & "/DDR_OUT",
            Xon            => Xon,
            MsgOn          => MsgOn,
            MsgSeverity    => WARNING);

          VitalSetupHoldCheck (
            Violation      => Tviol_DF_CLK_posedge,
            TimingData     => Tmkr_DF_CLK_posedge,
            TestSignal     => DF_ipd,
            TestSignalName => "DF",
            TestDelay      => 0 ns,
            RefSignal      => CLK_ipd,
            RefSignalName  => "CLK",
            RefDelay       => 0 ns,
            SetupHigh      => tsetup_DF_CLK_posedge_posedge,
            SetupLow       => tsetup_DF_CLK_negedge_posedge,
            HoldHigh       => thold_DF_CLK_posedge_posedge,
            HoldLow        => thold_DF_CLK_negedge_posedge,
            CheckEnabled   => TO_X01 (( NOT CLR_ipd )) /= '0',
            RefTransition  => 'R',
            HeaderMsg      => InstancePath & "/DDR_OUT",
            Xon            => Xon,
            MsgOn          => MsgOn,
            MsgSeverity    => WARNING);

          VitalRecoveryRemovalCheck (
            Violation      => Tviol_CLR_CLK_posedge,
            TimingData     => Tmkr_CLR_CLK_posedge,
            TestSignal     => CLR_ipd,
            TestSignalName => "CLR",
            TestDelay      => 0 ns,
            RefSignal      => CLK_ipd,
            RefSignalName  => "CLK",
            RefDelay       => 0 ns,
            Recovery       => trecovery_CLR_CLK_negedge_posedge,
            Removal        => thold_CLR_CLK_negedge_posedge,
            ActiveLow      => FALSE,
            CheckEnabled   => TRUE,
            RefTransition  => 'R',
            HeaderMsg      => InstancePath & "/DDR_OUT",
            Xon            => Xon,
            MsgOn          => MsgOn,
            MsgSeverity    => WARNING);

          VitalPeriodPulseCheck (
            Violation      => Pviol_CLK,
            PeriodData     => PInfo_CLK,
            TestSignal     => CLK_ipd,
            TestSignalName => "CLK",
            TestDelay      => 0 ns,
            Period         => tperiod_CLK_posedge,
            PulseWidthHigh => tpw_CLK_posedge,
            CheckEnabled   => TO_X01 ((( NOT CLR_ipd ))) /= '0',
            HeaderMsg      => InstancePath & "/DDR_OUT",
            Xon            => Xon,
            MsgOn          => MsgOn,
            MsgSeverity    => WARNING);

          VitalPeriodPulseCheck (
            Violation      => Pviol_CLR,
            PeriodData     => PInfo_CLR,
            TestSignal     => CLR_ipd,
            TestSignalName => "CLR",
            TestDelay      => 0 ns,
            Period         => 0 ns,
            PulseWidthHigh => tpw_CLR_posedge,
            PulseWidthLow  => 0 ns,
            CheckEnabled   => TRUE,
            HeaderMsg      => InstancePath & "/DDR_OUT",
            Xon            => Xon,
            MsgOn          => MsgOn,
            MsgSeverity    => WARNING);

        end if;

        --------------------------------
        --  Functionality Section
        -------------------------------

        Violation := Tviol_DR_CLK_posedge or Tviol_DF_CLK_posedge or Tviol_CLR_CLK_posedge;

        VitalStateTable(
          Result => QR_tmp,
          PreviousDataIn => PrevData_QR,
          StateTable => DFN1C1_Q_tab,
          DataIn => ( CLR_ipd, CLK_ipd, DR_ipd ));
        QR_tmp := Violation XOR QR_tmp;

        VitalStateTable(
          Result => QF_tmp,
          PreviousDataIn => PrevData_QF,
          StateTable => DFN1C1_Q_tab,
          DataIn => ( CLR_ipd, CLK_ipd, DF_ipd ));
        QF_tmp := Violation XOR QF_tmp;

        Q_zd := VitalMUX2( QR_tmp, QF_tmp, CLK_ipd );

        ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
          OutSignal     => Q,
          GlitchData    => Q_GlitchData,
          OutSignalName => "Q",
          OutTemp       => Q_zd,
          Paths         => ( 0 => ( CLK_ipd'last_event, tpd_CLK_Q, true ),
                             1 => ( CLR_ipd'last_event, tpd_CLR_Q, true )),
          Mode          => OnDetect,
          Xon           => Xon,
          MsgOn         => MsgOn,
          MsgSeverity   => WARNING);

  end process;

end VITAL_ACT;

configuration CFG_DDR_OUT_VITAL of DDR_OUT is
  for VITAL_ACT
  end for;
end CFG_DDR_OUT_VITAL;

 ---- CELL DDR_REG ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DDR_REG is
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_QR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_QF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLK_QR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLK_QF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tsetup_D_CLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_D_CLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_D_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_D_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_CLR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_CLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_CLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_D        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));

 
  port(
                CLR             :   in    STD_ULOGIC;
                CLK            :   in    STD_ULOGIC;
                D             :  in    STD_ULOGIC;
                QF               :  out    STD_ULOGIC;
                QR               :  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DDR_REG :  entity is TRUE;
 end DDR_REG;




-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of DDR_REG is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL D_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
          VitalWireDelay (D_ipd, D, tipd_D);
          VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
          VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
        end block;



  --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

        -- timing check results
        VARIABLE Tviol_D_CLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_D_CLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_CLR_CLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_CLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Pviol_CLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_CLK     : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_CLR      : STD_ULOGIC := '0';
        VARIABLE PInfo_CLR      : VitalPeriodDataType := VitalPeriodDataInit;

        -- functionality results
        VARIABLE Violation      : STD_ULOGIC := '0';
        VARIABLE PrevData_Qtmp  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 6);

        VARIABLE CLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE D_delayed    : STD_ULOGIC := 'X';
        VARIABLE tmp_zd    : STD_ULOGIC := 'X';

        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');

        ALIAS QR_zd : STD_LOGIC is Results(1);
        ALIAS QF_zd : STD_LOGIC is Results(2);


        -- output glitch detection variables
        VARIABLE QR_GlitchData  : VitalGlitchDataType;
        VARIABLE QF_GlitchData  : VitalGlitchDataType;

   begin
  ------------------------
   --  Timing Check Section
   ------------------------

  if(TimingChecksOn) then
        VitalSetupHoldCheck (
         Violation              => Tviol_D_CLK_posedge,
         TimingData             => Tmkr_D_CLK_posedge,
         TestSignal             => D_ipd,
         TestSignalName         => "D",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_D_CLK_posedge_posedge,
         SetupLow               => tsetup_D_CLK_negedge_posedge,
         HoldHigh               => thold_D_CLK_posedge_posedge,
         HoldLow                => thold_D_CLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/DDR_REG",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);



        VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_CLK_posedge,
         TimingData             => Tmkr_CLR_CLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_CLK_negedge_posedge,
         Removal               => thold_CLR_CLK_negedge_posedge,
         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "DDR_REG",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


        VitalPeriodPulseCheck (
         Violation              => Pviol_CLK,
         PeriodData             => PInfo_CLK,
         TestSignal             => CLK_ipd,
         TestSignalName         => "CLK",
         TestDelay              => 0 ns,
         Period         => tperiod_CLK_posedge,
         PulseWidthLow  => tpw_CLK_negedge,
         PulseWidthHigh => tpw_CLK_posedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "DDR_REG",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


       VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period         => 0 ns,
         PulseWidthHigh => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "DDR_REG",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        end if;


      --------------------------------
      --  Functionality Section
      -------------------------------


      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge;

      VitalStateTable(
       Result => tmp_zd,
       PreviousDataIn => PrevData_Qtmp,
       StateTable => DFEG_Q_tab,
       DataIn => (
             '1', CLK_ipd, tmp_zd, D_delayed,  '0', '1', CLK_delayed));
       tmp_zd := Violation XOR tmp_zd;

      VitalStateTable(
       Result => QF_zd,
       PreviousDataIn => PrevData_QF,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), CLK_delayed, QF_zd, tmp_zd, '0', '1', CLK_ipd));
       QF_zd := Violation XOR QF_zd;

       VitalStateTable(
       Result => QR_zd,
       PreviousDataIn => PrevData_QR,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), CLK_delayed, QR_zd, D_delayed, '0', '1', CLK_ipd));
       QR_zd := Violation XOR QR_zd;

       D_delayed := D_ipd;
       CLK_delayed := CLK_ipd;


        ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
         OutSignal => QR,
         GlitchData => QR_GlitchData,
         OutSignalName => "QR",
         OutTemp => QR_zd,
         Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QR, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_QR, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

       VitalPathDelay01 (
         OutSignal => QF,
         GlitchData => QF_GlitchData,
         OutSignalName => "QF",
         OutTemp => QF_zd,
         Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QF, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_QF, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

 end process;


end VITAL_ACT;

configuration CFG_DDR_REG_VITAL of DDR_REG is
   for VITAL_ACT
   end for;
end CFG_DDR_REG_VITAL;


---- CELL IOBI_ID_OB_EB ----
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
 entity IOBI_ID_OB_EB is
   generic (
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;

      tipd_D           : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E           : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ICLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_YIN         : VitalDelayType01 := (0.000 ns, 0.000 ns);

      tpd_D_DOUT       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_E_EOUT       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLR_YR       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLR_YF       : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_ICLK_YR      : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_ICLK_YF      : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_YIN_ICLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_YIN_ICLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_negedge_posedge     : VitalDelayType := 0.000 ns;

      tsetup_YIN_ICLK_posedge_negedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_posedge_negedge     : VitalDelayType := 0.000 ns;
      tsetup_YIN_ICLK_negedge_negedge    : VitalDelayType := 0.000 ns;
      thold_YIN_ICLK_negedge_negedge     : VitalDelayType := 0.000 ns;

      trecovery_CLR_ICLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_CLR_ICLK_negedge_posedge     : VitalDelayType := 0.000 ns;

      tpw_ICLK_posedge                   :  VitalDelayType := 0.000 ns;
      tpw_ICLK_negedge                   :  VitalDelayType := 0.000 ns;
      tperiod_ICLK_posedge               :  VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                    :  VitalDelayType := 0.000 ns
     );


   port (
      D             :  in    std_ulogic;
      CLR           :  in    std_ulogic;
      E             :  in    std_ulogic;
      ICLK          :  in    std_ulogic;
      YIN           :  in    std_ulogic;
      DOUT          :  out   std_ulogic;
      EOUT          :  out   std_ulogic;
      YR            :  out   std_ulogic;
      YF            :  out   std_ulogic
     );

   attribute VITAL_LEVEL0 of IOBI_ID_OB_EB :  entity is TRUE;
   
end IOBI_ID_OB_EB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_ID_OB_EB is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

  signal D_ipd    : std_ulogic := 'X';
  signal CLR_ipd  : std_ulogic := 'X';
  signal E_ipd    : std_ulogic := 'X';
  signal ICLK_ipd : std_ulogic := 'X';
  signal YIN_ipd  : std_ulogic := 'X';

  begin  --  VITAL_ACT
  
  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WireDelay: block

  begin  --  block WireDelay
  
    VitalWireDelay (D_ipd,    D,    VitalExtendToFillDelay(tipd_D));
    VitalWireDelay (CLR_ipd,  CLR,  VitalExtendToFillDelay(tipd_CLR));
    VitalWireDelay (E_ipd,    E,    VitalExtendToFillDelay(tipd_E));
    VitalWireDelay (ICLK_ipd, ICLK, VitalExtendToFillDelay(tipd_ICLK));
    VitalWireDelay (YIN_ipd,  YIN,  VitalExtendToFillDelay(tipd_YIN));
    
  end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################
  VITALBehavior : process (D_ipd, CLR_ipd, E_ipd, ICLK_ipd, YIN_ipd)


    -- timing check results
    variable Tviol_YIN_ICLK_posedge : std_ulogic := '0';
    variable Tmkr_YIN_ICLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
    variable Tviol_YIN_ICLK_negedge : std_ulogic := '0';
    variable Tmkr_YIN_ICLK_negedge  : VitalTimingDataType := VitalTimingDataInit;
    variable Tviol_CLR_ICLK_posedge : std_ulogic := '0';
    variable Tmkr_CLR_ICLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
    variable Pviol_ICLK             : std_ulogic := '0';
    variable PInfo_ICLK             : VitalPeriodDataType := VitalPeriodDataInit;
    variable Pviol_CLR              : std_ulogic := '0';
    variable PInfo_CLR              : VitalPeriodDataType := VitalPeriodDataInit;

    -- functionality results
    variable Violation              : std_ulogic := '0';
    variable PrevData_Qtmp          : STD_LOGIC_VECTOR(0 to 6);
    variable PrevData_QR            : STD_LOGIC_VECTOR(0 to 6);
    variable PrevData_QF            : STD_LOGIC_VECTOR(0 to 6);

    variable ICLK_delayed           : std_ulogic := 'X';
    variable YIN_delayed            : std_ulogic := 'X';

    variable DOUT_zd                : std_ulogic := 'X';
    variable EOUT_zd                : std_ulogic := 'X';
    variable tmp_zd                 : std_ulogic := 'X';
    variable YR_zd                  : std_ulogic := 'X';
    variable YF_zd                  : std_ulogic := 'X';

    -- output glitch detection variables
    variable DOUT_GlitchData        : VitalGlitchDataType;
    variable EOUT_GlitchData        : VitalGlitchDataType;
    variable YR_GlitchData          : VitalGlitchDataType;
    variable YF_GlitchData          : VitalGlitchDataType;


  begin

  
    ------------------------
    --  Timing Check Section
    ------------------------

    if (TimingChecksOn) then
       VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_posedge,
         TimingData             => Tmkr_YIN_ICLK_posedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
         HoldHigh               => thold_YIN_ICLK_posedge_posedge,
         HoldLow                => thold_YIN_ICLK_negedge_posedge,
         CheckEnabled           => TO_X01(CLR_ipd) /= '1',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OB_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_negedge,
         TimingData             => Tmkr_YIN_ICLK_negedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_negedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_negedge,
         HoldHigh               => thold_YIN_ICLK_posedge_negedge,
         HoldLow                => thold_YIN_ICLK_negedge_negedge,
         CheckEnabled           => TO_X01(CLR_ipd) /= '1',
         RefTransition          => 'F',
         HeaderMsg              => InstancePath & "/IOBI_ID_OB_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

       VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_ICLK_posedge,
         TimingData             => Tmkr_CLR_ICLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         Recovery               => trecovery_CLR_ICLK_negedge_posedge,
         Removal                => thold_CLR_ICLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "IOBI_ID_OB_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

       VitalPeriodPulseCheck (
         Violation              => Pviol_ICLK,
         PeriodData             => PInfo_ICLK,
         TestSignal             => ICLK_ipd,
         TestSignalName         => "ICLK",
         TestDelay              => 0 ns,
         Period                 => tperiod_ICLK_posedge,
         PulseWidthHigh         => tpw_ICLK_posedge,
         PulseWidthLow          => tpw_ICLK_negedge,
         CheckEnabled           => TO_X01(CLR_ipd) /= '1',
         HeaderMsg              => InstancePath & "IOBI_ID_OB_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);


       VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period                 => 0 ns,
         PulseWidthHigh         => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOBI_ID_OB_EB",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

    end if;
    
    --------------------------------
    --  Functionality Section
    -------------------------------

    Violation := Tviol_YIN_ICLK_posedge or Tviol_YIN_ICLK_negedge or 
                 Tviol_CLR_ICLK_posedge or Pviol_ICLK or Pviol_CLR;

    DOUT_zd := TO_X01(D_ipd);
    EOUT_zd := TO_X01(E_ipd);

    VitalStateTable(
      Result => tmp_zd,
      PreviousDataIn => PrevData_Qtmp,
      StateTable => DFEG_Q_tab,
      DataIn => (
             '1', (NOT ICLK_delayed), tmp_zd, YIN_delayed, '0', '1', (NOT ICLK_ipd)));
      tmp_zd := Violation XOR tmp_zd;

    VitalStateTable(
      Result => YF_zd,
      PreviousDataIn => PrevData_QF,
      StateTable => DFEG_Q_tab,
      DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YF_zd, tmp_zd, '0', '1', ICLK_ipd));
      YF_zd := Violation XOR YF_zd;

    VitalStateTable(
      Result => YR_zd,
      PreviousDataIn => PrevData_QR,
      StateTable => DFEG_Q_tab,
      DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YR_zd, YIN_delayed, '0', '1', ICLK_ipd));
      YR_zd := Violation XOR YR_zd;

    ICLK_delayed := ICLK_ipd;
    YIN_delayed  := YIN_ipd;
    
    ----------------------
    --  Path Delay Section
    ----------------------
    
    VitalPathDelay01 (
         OutSignal     => DOUT,
         GlitchData    => DOUT_GlitchData,
         OutSignalName => "DOUT",
         OutTemp       => DOUT_zd,
         Paths         => (0 => (D_ipd'last_event, tpd_D_DOUT, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

    VitalPathDelay01 (
         OutSignal     => EOUT,
         GlitchData    => EOUT_GlitchData,
         OutSignalName => "EOUT",
         OutTemp       => EOUT_zd,
         Paths         => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

    VitalPathDelay01 (
         OutSignal     => YR,
         GlitchData    => YR_GlitchData,
         OutSignalName => "YR",
         OutTemp       => YR_zd,
         Paths         => (0 => (ICLK_ipd'last_event, tpd_ICLK_YR, true),
                           1 => (CLR_ipd'last_event,  tpd_CLR_YR,  true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

    VitalPathDelay01 (
         OutSignal     => YF,
         GlitchData    => YF_GlitchData,
         OutSignalName => "YF",
         OutTemp       => YF_zd,
         Paths         => (0 => (ICLK_ipd'last_event, tpd_ICLK_YF, true),
                           1 => (CLR_ipd'last_event,  tpd_CLR_YF,  true)),
         Mode          => OnDetect,
         Xon           => Xon,
         MsgOn         => MsgOn,
         MsgSeverity   => WARNING);

  end process;

end VITAL_ACT;

configuration CFG_IOBI_ID_OB_EB_VITAL of IOBI_ID_OB_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_ID_OB_EB_VITAL;


---- CELL IOBI_ID_OD_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_ID_OD_EB is
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_EOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_YIN_ICLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_YIN_ICLK_posedge_negedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;



                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                thold_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_ICLK_posedge    :  VitalDelayType := 0.000 ns;

                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;

                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_YIN        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_ICLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                ICLK            :   in    STD_ULOGIC;
                YIN             :   in    STD_ULOGIC;
                E               :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                YR               :  out    STD_ULOGIC;
                YF               :  out    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOBI_ID_OD_EB :  entity is TRUE;
 end IOBI_ID_OD_EB;

 -- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_ID_OD_EB is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL DR_ipd  : STD_ULOGIC := 'X';
        SIGNAL DF_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
        SIGNAL OCLK_ipd : STD_ULOGIC := 'X';
        SIGNAL ICLK_ipd : STD_ULOGIC := 'X';


  begin

               ---------------------
               --  INPUT PATH DELAYs
               ---------------------
               WireDelay : block
               begin
                 VitalWireDelay (DR_ipd, DR, tipd_DR);
                 VitalWireDelay (DF_ipd, DF, tipd_DF);
                 VitalWireDelay (E_ipd, E, tipd_E);
                 VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
                 VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
                 VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
                 VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
               end block;

    --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (DR_ipd, DF_ipd,YIN_ipd,E_ipd,CLR_ipd,ICLK_ipd, OCLK_ipd)


        -- timing check results
        VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_YIN_ICLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_YIN_ICLK_negedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_YIN_ICLK_negedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_DR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_DF_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DF_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_ICLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Pviol_OCLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_OCLK     : VitalPeriodDataType := VitalPeriodDataInit;

        VARIABLE Pviol_ICLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_ICLK     : VitalPeriodDataType := VitalPeriodDataInit;

        VARIABLE Pviol_CLR      : STD_ULOGIC := '0';
        VARIABLE PInfo_CLR      : VitalPeriodDataType := VitalPeriodDataInit;

        -- functionality results
        VARIABLE Violation      : STD_ULOGIC := '0';
        VARIABLE PrevData_Qtmp  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE PrevData_QR2  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QF2  : STD_LOGIC_VECTOR(0 to 6);

        VARIABLE OCLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE ICLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE YIN_delayed    : STD_ULOGIC := 'X';


        VARIABLE E_delayed    : STD_ULOGIC := 'X';

        VARIABLE DR_tmp    : STD_ULOGIC := 'X';
        VARIABLE DF_tmp    : STD_ULOGIC := 'X';
        VARIABLE tmp_zd    : STD_ULOGIC := 'X';

        VARIABLE Results : STD_LOGIC_VECTOR(1 to 4)  := (others => 'X');

        ALIAS DOUT_zd : STD_LOGIC is Results(1);
        ALIAS YR_zd : STD_LOGIC is Results(2);
        ALIAS YF_zd : STD_LOGIC is Results(3);
        ALIAS EOUT_zd : STD_LOGIC is Results(4);

        -- output glitch detection variables
        VARIABLE YR_GlitchData  : VitalGlitchDataType;
        VARIABLE YF_GlitchData  : VitalGlitchDataType;
        VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
        VARIABLE EOUT_GlitchData  : VitalGlitchDataType;


   begin

  
   ------------------------
   --  Timing Check Section
   ------------------------

   if(TimingChecksOn) then
        VitalSetupHoldCheck (
         Violation              => Tviol_DR_OCLK_posedge,
         TimingData             => Tmkr_DR_OCLK_posedge,
         TestSignal             => DR_ipd,
         TestSignalName         => "DR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DR_OCLK_posedge_posedge,
         SetupLow               => tsetup_DR_OCLK_negedge_posedge,
         HoldHigh               => thold_DR_OCLK_posedge_posedge,
         HoldLow                => thold_DR_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


         VitalSetupHoldCheck (
         Violation              => Tviol_DF_OCLK_posedge,
         TimingData             => Tmkr_DF_OCLK_posedge,
         TestSignal             => DF_ipd,
         TestSignalName         => "DF",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DF_OCLK_posedge_posedge,
         SetupLow               => tsetup_DF_OCLK_negedge_posedge,
         HoldHigh               => thold_DF_OCLK_posedge_posedge,
         HoldLow                => thold_DF_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_posedge,
         TimingData             => Tmkr_YIN_ICLK_posedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
         HoldHigh               => thold_YIN_ICLK_posedge_posedge,
         HoldLow                => thold_YIN_ICLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);



         VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_negedge,
         TimingData             => Tmkr_YIN_ICLK_negedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_negedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_negedge,
         HoldHigh               => thold_YIN_ICLK_posedge_negedge,
         HoldLow                => thold_YIN_ICLK_negedge_negedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'F',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


        VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_OCLK_posedge,
         TimingData             => Tmkr_CLR_OCLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_OCLK_negedge_posedge,
         Removal               => thold_CLR_OCLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

       VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_ICLK_posedge,
         TimingData             => Tmkr_CLR_ICLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_ICLK_negedge_posedge,
         Removal               => thold_CLR_ICLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


        VitalPeriodPulseCheck (
         Violation              => Pviol_OCLK,
         PeriodData             => PInfo_OCLK,
         TestSignal             => OCLK_ipd,
         TestSignalName         => "OCLK",
         TestDelay              => 0 ns,
         Period         => tperiod_OCLK_posedge,
         PulseWidthHigh => tpw_OCLK_posedge,
         PulseWidthLow  => tpw_OCLK_negedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


       VitalPeriodPulseCheck (
         Violation              => Pviol_ICLK,
         PeriodData             => PInfo_ICLK,
         TestSignal             => ICLK_ipd,
         TestSignalName         => "ICLK",
         TestDelay              => 0 ns,
         Period         => tperiod_ICLK_posedge,
         PulseWidthHigh => tpw_ICLK_posedge,
         PulseWidthLow  => tpw_ICLK_negedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


         VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period         => 0 ns,
         PulseWidthHigh => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        end if;

  

      --------------------------------
      --  Functionality Section
      -------------------------------

   Violation := Tviol_DR_OCLK_posedge or Tviol_DF_OCLK_posedge or Tviol_CLR_OCLK_posedge or Tviol_YIN_ICLK_posedge or Tviol_CLR_ICLK_posedge;

      VitalStateTable(
       Result => DR_tmp,
       PreviousDataIn => PrevData_QR,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DR_ipd ));
       DR_tmp := Violation XOR DR_tmp;

      VitalStateTable(
       Result => DF_tmp,
       PreviousDataIn => PrevData_QF,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DF_ipd ));
       DF_tmp := Violation XOR DF_tmp;

      DOUT_zd := VitalMUX2( DR_tmp, DF_tmp, OCLK_ipd );
      EOUT_zd :=TO_X01(E_delayed);




      VitalStateTable(
       Result => tmp_zd,
       PreviousDataIn => PrevData_Qtmp,
       StateTable => DFEG_Q_tab,
       DataIn => (
             '1', ICLK_ipd, tmp_zd, YIN_delayed,  '0', '1', ICLK_delayed));
       tmp_zd := Violation XOR tmp_zd;

      VitalStateTable(
       Result => YF_zd,
       PreviousDataIn => PrevData_QF2,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YF_zd, tmp_zd, '0', '1', ICLK_ipd));
       YF_zd := Violation XOR YF_zd;

       VitalStateTable(
       Result => YR_zd,
       PreviousDataIn => PrevData_QR2,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YR_zd, YIN_delayed, '0', '1', ICLK_ipd));
       YR_zd := Violation XOR YR_zd;

      YIN_delayed := YIN_ipd;
      ICLK_delayed := ICLK_ipd;
      E_delayed  := E_ipd;
      OCLK_delayed :=OCLK_ipd;



       ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
         OutSignal => DOUT,
         GlitchData => DOUT_GlitchData,
         OutSignalName => "DOUT",
         OutTemp => DOUT_zd,
         Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

       VitalPathDelay01 (
         OutSignal => EOUT,
         GlitchData => EOUT_GlitchData,
         OutSignalName => "EOUT",
         OutTemp => EOUT_zd,
         Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

        VitalPathDelay01 (
         OutSignal => YR,
         GlitchData => YR_GlitchData,
         OutSignalName => "YR",
         OutTemp => YR_zd,
         Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_YR, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_YR, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

  VitalPathDelay01 (
         OutSignal => YF,
         GlitchData => YF_GlitchData,
         OutSignalName => "YF",
         OutTemp => YF_zd,
         Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_YF, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_YF, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);



   end process;

end VITAL_ACT;

configuration CFG_IOBI_ID_OD_EB_VITAL of IOBI_ID_OD_EB is
   for VITAL_ACT
   end for;
end CFG_IOBI_ID_OD_EB_VITAL;



---- CELL IOBI_ID_OD_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBI_ID_OD_ERC is
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_EOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_EOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tpd_CLR_YR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_YIN_ICLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_YIN_ICLK_posedge_negedge :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_E_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;



                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                thold_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_ICLK_posedge    :  VitalDelayType := 0.000 ns;

                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge    :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_YIN        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_ICLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                ICLK            :   in    STD_ULOGIC;
                YIN             :   in    STD_ULOGIC;
                E               :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                YR               :  out    STD_ULOGIC;
                YF               :  out    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOBI_ID_OD_ERC :  entity is TRUE;
 end IOBI_ID_OD_ERC;

 -- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOBI_ID_OD_ERC is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL DR_ipd  : STD_ULOGIC := 'X';
        SIGNAL DF_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
        SIGNAL OCLK_ipd : STD_ULOGIC := 'X';
        SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

   begin

               ---------------------
                 --  INPUT PATH DELAYs
                 ---------------------
                 WireDelay : block
                 begin
                   VitalWireDelay (DR_ipd, DR, tipd_DR);
                   VitalWireDelay (DF_ipd, DF, tipd_DF);
                   VitalWireDelay (E_ipd, E, tipd_E);
                   VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
                   VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
                   VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
                   VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
                 end block;



   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (DR_ipd, DF_ipd,YIN_ipd,E_ipd,CLR_ipd,ICLK_ipd, OCLK_ipd)

        -- timing check results
        VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_YIN_ICLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_YIN_ICLK_negedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_YIN_ICLK_negedge : VitalTimingDataType := VitalTimingDataInit;


        VARIABLE Tviol_DR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_DF_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DF_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_E_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_ICLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Pviol_OCLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_OCLK     : VitalPeriodDataType := VitalPeriodDataInit;

        VARIABLE Pviol_ICLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_ICLK     : VitalPeriodDataType := VitalPeriodDataInit;

        VARIABLE Pviol_CLR      : STD_ULOGIC := '0';
        VARIABLE PInfo_CLR      : VitalPeriodDataType := VitalPeriodDataInit;

        -- functionality results
        VARIABLE Violation      : STD_ULOGIC := '0';
        VARIABLE PrevData_Qtmp  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE PrevData_QR2  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QF2  : STD_LOGIC_VECTOR(0 to 6);

        VARIABLE PrevData_QE  : STD_LOGIC_VECTOR(0 to 6);

        VARIABLE OCLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE ICLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE YIN_delayed    : STD_ULOGIC := 'X';

        VARIABLE E_delayed    : STD_ULOGIC := 'X';

        VARIABLE DR_tmp    : STD_ULOGIC := 'X';
        VARIABLE DF_tmp    : STD_ULOGIC := 'X';
        VARIABLE tmp_zd    : STD_ULOGIC := 'X';

        VARIABLE Results : STD_LOGIC_VECTOR(1 to 4)  := (others => 'X');

        ALIAS DOUT_zd : STD_LOGIC is Results(1);
        ALIAS YR_zd : STD_LOGIC is Results(2);
        ALIAS YF_zd : STD_LOGIC is Results(3);
        ALIAS EOUT_zd : STD_LOGIC is Results(4);

        -- output glitch detection variables
        VARIABLE YR_GlitchData  : VitalGlitchDataType;
        VARIABLE YF_GlitchData  : VitalGlitchDataType;
        VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
        VARIABLE EOUT_GlitchData  : VitalGlitchDataType;


   begin

 ------------------------
   --  Timing Check Section
   ------------------------

   if(TimingChecksOn) then
        VitalSetupHoldCheck (
         Violation              => Tviol_DR_OCLK_posedge,
         TimingData             => Tmkr_DR_OCLK_posedge,
         TestSignal             => DR_ipd,
         TestSignalName         => "DR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DR_OCLK_posedge_posedge,
         SetupLow               => tsetup_DR_OCLK_negedge_posedge,
         HoldHigh               => thold_DR_OCLK_posedge_posedge,
         HoldLow                => thold_DR_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


       VitalSetupHoldCheck (
         Violation              => Tviol_DF_OCLK_posedge,
         TimingData             => Tmkr_DF_OCLK_posedge,
         TestSignal             => DF_ipd,
         TestSignalName         => "DF",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DF_OCLK_posedge_posedge,
         SetupLow               => tsetup_DF_OCLK_negedge_posedge,
         HoldHigh               => thold_DF_OCLK_posedge_posedge,
         HoldLow                => thold_DF_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


       VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_posedge,
         TimingData             => Tmkr_YIN_ICLK_posedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
         HoldHigh               => thold_YIN_ICLK_posedge_posedge,
         HoldLow                => thold_YIN_ICLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


       VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_negedge,
         TimingData             => Tmkr_YIN_ICLK_negedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_negedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_negedge,
         HoldHigh               => thold_YIN_ICLK_posedge_negedge,
         HoldLow                => thold_YIN_ICLK_negedge_negedge,
         CheckEnabled           =>
         TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'F',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);




       VitalSetupHoldCheck (
         Violation              => Tviol_E_OCLK_posedge,
         TimingData             => Tmkr_E_OCLK_posedge,
         TestSignal             => E_ipd,
         TestSignalName         => "E",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_E_OCLK_posedge_posedge,
         SetupLow               => tsetup_E_OCLK_negedge_posedge,
         HoldHigh               => thold_E_OCLK_posedge_posedge,
         HoldLow                => thold_E_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


        VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_OCLK_posedge,
         TimingData             => Tmkr_CLR_OCLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_OCLK_negedge_posedge,
         Removal               => thold_CLR_OCLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

       VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_ICLK_posedge,
         TimingData             => Tmkr_CLR_ICLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_ICLK_negedge_posedge,
         Removal               => thold_CLR_ICLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);



         VitalPeriodPulseCheck (
         Violation              => Pviol_ICLK,
         PeriodData             => PInfo_ICLK,
         TestSignal             => ICLK_ipd,
         TestSignalName         => "ICLK",
         TestDelay              => 0 ns,
         Period         => tperiod_ICLK_posedge,
         PulseWidthHigh => tpw_ICLK_posedge,
         PulseWidthLow  => tpw_ICLK_negedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        VitalPeriodPulseCheck (
          Violation              => Pviol_OCLK,
          PeriodData             => PInfo_OCLK,
          TestSignal             => OCLK_ipd,
          TestSignalName         => "OCLK",
          TestDelay              => 0 ns,
          Period         => tperiod_OCLK_posedge,
          PulseWidthHigh => tpw_OCLK_posedge,
          PulseWidthLow  => tpw_OCLK_negedge,
          CheckEnabled           =>
          TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
          Xon            => Xon,
          MsgOn          => MsgOn,
          MsgSeverity            => WARNING);

         

         VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period         => 0 ns,
         PulseWidthHigh => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOBI_ID_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        end if;
      --------------------------------
      --  Functionality Section
      -------------------------------

    Violation := Tviol_DR_OCLK_posedge or Tviol_DF_OCLK_posedge or Tviol_CLR_OCLK_posedge or Tviol_YIN_ICLK_posedge or Tviol_CLR_ICLK_posedge or Tviol_E_OCLK_posedge;

      VitalStateTable(
       Result => DR_tmp,
       PreviousDataIn => PrevData_QR,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DR_ipd ));
       DR_tmp := Violation XOR DR_tmp;

      VitalStateTable(
       Result => DF_tmp,
       PreviousDataIn => PrevData_QF,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DF_ipd ));
       DF_tmp := Violation XOR DF_tmp;

      DOUT_zd := VitalMUX2( DR_tmp, DF_tmp, OCLK_ipd );

      VitalStateTable(
       Result => EOUT_zd,
       PreviousDataIn => PrevData_QE,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  '0', '1', ICLK_ipd));
       EOUT_zd := Violation XOR EOUT_zd;

      VitalStateTable(
       Result => tmp_zd,
       PreviousDataIn => PrevData_Qtmp,
       StateTable => DFEG_Q_tab,
       DataIn => (
             '1', ICLK_ipd, tmp_zd, YIN_delayed,  '0', '1', ICLK_delayed));
       tmp_zd := Violation XOR tmp_zd;

      VitalStateTable(
       Result => YF_zd,
       PreviousDataIn => PrevData_QF2,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YF_zd, tmp_zd, '0', '1', ICLK_ipd));
       YF_zd := Violation XOR YF_zd;

       VitalStateTable(
       Result => YR_zd,
       PreviousDataIn => PrevData_QR2,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YR_zd, YIN_delayed, '0', '1', ICLK_ipd));
       YR_zd := Violation XOR YR_zd;

      YIN_delayed := YIN_ipd;
      ICLK_delayed := ICLK_ipd;
      E_delayed  := E_ipd;
      OCLK_delayed :=OCLK_ipd;


   
  
       ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
         OutSignal => DOUT,
         GlitchData => DOUT_GlitchData,
         OutSignalName => "DOUT",
         OutTemp => DOUT_zd,
         Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

       VitalPathDelay01 (
         OutSignal => EOUT,
         GlitchData => EOUT_GlitchData,
         OutSignalName => "EOUT",
         OutTemp => EOUT_zd,
         Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_EOUT, true)),

         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

        VitalPathDelay01 (
         OutSignal => YR,
         GlitchData => YR_GlitchData,
         OutSignalName => "YR",
         OutTemp => YR_zd,
         Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_YR, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_YR, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);
    VitalPathDelay01 (
         OutSignal => YF,
         GlitchData => YF_GlitchData,
         OutSignalName => "YF",
         OutTemp => YF_zd,
         Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_YF, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_YF, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);



   end process;

end VITAL_ACT;

configuration CFG_IOBI_ID_OD_ERC_VITAL of IOBI_ID_OD_ERC is
   for VITAL_ACT
   end for;
end CFG_IOBI_ID_OD_ERC_VITAL;

 ---- CELL IOIN_ID ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOIN_ID is
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_YR      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_YF      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YR     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_ICLK_YF     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_YIN_ICLK_posedge_posedge  :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_posedge  :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_posedge_negedge  :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_posedge_negedge   :   VitalDelayType := 0.000 ns;
                tsetup_YIN_ICLK_negedge_negedge  :   VitalDelayType := 0.000 ns;
                thold_YIN_ICLK_negedge_negedge   :   VitalDelayType := 0.000 ns;

                thold_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_ICLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_ICLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_ICLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_ICLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_YIN        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_ICLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));

  
  port(
                CLR             :   in    STD_ULOGIC;
                ICLK            :   in    STD_ULOGIC;
                YIN             :  in    STD_ULOGIC;
                YF               :  out    STD_ULOGIC;
                YR               :  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOIN_ID :  entity is TRUE;
 end IOIN_ID;



-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOIN_ID is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL YIN_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
        SIGNAL ICLK_ipd : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
          VitalWireDelay (YIN_ipd, YIN, tipd_YIN);
          VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
          VitalWireDelay (ICLK_ipd,ICLK, tipd_ICLK);
        end block;


  --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (YIN_ipd, CLR_ipd,ICLK_ipd)

        -- timing check results
        VARIABLE Tviol_YIN_ICLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_YIN_ICLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_YIN_ICLK_negedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_YIN_ICLK_negedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_CLR_ICLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_ICLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Pviol_ICLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_ICLK     : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_CLR      : STD_ULOGIC := '0';
        VARIABLE PInfo_CLR      : VitalPeriodDataType := VitalPeriodDataInit;

        -- functionality results
        VARIABLE Violation      : STD_ULOGIC := '0';
        VARIABLE PrevData_Qtmp  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 6);

        VARIABLE ICLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE YIN_delayed    : STD_ULOGIC := 'X';
        VARIABLE tmp_zd    : STD_ULOGIC := 'X';

        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');

        ALIAS YR_zd : STD_LOGIC is Results(1);
        ALIAS YF_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE YR_GlitchData  : VitalGlitchDataType;
        VARIABLE YF_GlitchData  : VitalGlitchDataType;

   begin

  ------------------------
   --  Timing Check Section
   ------------------------

  if(TimingChecksOn) then
        VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_posedge,
         TimingData             => Tmkr_YIN_ICLK_posedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_posedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_posedge,
         HoldHigh               => thold_YIN_ICLK_posedge_posedge,
         HoldLow                => thold_YIN_ICLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOIN_ID",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

        VitalSetupHoldCheck (
         Violation              => Tviol_YIN_ICLK_negedge,
         TimingData             => Tmkr_YIN_ICLK_negedge,
         TestSignal             => YIN_ipd,
         TestSignalName         => "YIN",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_YIN_ICLK_posedge_negedge,
         SetupLow               => tsetup_YIN_ICLK_negedge_negedge,
         HoldHigh               => thold_YIN_ICLK_posedge_negedge,
         HoldLow                => thold_YIN_ICLK_negedge_negedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'F',
         HeaderMsg              => InstancePath & "/IOIN_ID",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


        VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_ICLK_posedge,
         TimingData             => Tmkr_CLR_ICLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => ICLK_ipd,
         RefSignalName          => "ICLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_ICLK_negedge_posedge,
         Removal               => thold_CLR_ICLK_negedge_posedge,
         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOIN_ID",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        VitalPeriodPulseCheck (
         Violation              => Pviol_ICLK,
         PeriodData             => PInfo_ICLK,
         TestSignal             => ICLK_ipd,
         TestSignalName         => "ICLK",
         TestDelay              => 0 ns,
         Period         => tperiod_ICLK_posedge,
         PulseWidthHigh => tpw_ICLK_posedge,
         PulseWidthLow  => tpw_ICLK_negedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOIN_ID",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


       VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period         => 0 ns,
         PulseWidthHigh => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOIN_ID",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        end if;


      --------------------------------
      --  Functionality Section
      -------------------------------

        Violation := Tviol_YIN_ICLK_posedge or Tviol_CLR_ICLK_posedge;

      VitalStateTable(
       Result => tmp_zd,
       PreviousDataIn => PrevData_Qtmp,
       StateTable => DFEG_Q_tab,
       DataIn => (
             '1', ICLK_ipd, tmp_zd, YIN_delayed,  '0', '1', ICLK_delayed));
       tmp_zd := Violation XOR tmp_zd;

      VitalStateTable(
       Result => YF_zd,
       PreviousDataIn => PrevData_QF,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YF_zd, tmp_zd, '0', '1', ICLK_ipd));
       YF_zd := Violation XOR YF_zd;

       VitalStateTable(
       Result => YR_zd,
       PreviousDataIn => PrevData_QR,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), ICLK_delayed, YR_zd, YIN_delayed, '0', '1', ICLK_ipd));
       YR_zd := Violation XOR YR_zd;

     YIN_delayed := YIN_ipd;
     ICLK_delayed := ICLK_ipd;



       ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
         OutSignal => YR,
         GlitchData => YR_GlitchData,
         OutSignalName => "YR",
         OutTemp => YR_zd,
         Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_YR, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_YR, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

       VitalPathDelay01 (
         OutSignal => YF,
         GlitchData => YF_GlitchData,
         OutSignalName => "YF",
         OutTemp => YF_zd,
         Paths => (0 => (ICLK_ipd'last_event, tpd_ICLK_YF, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_YF, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOIN_ID_VITAL of IOIN_ID is
   for VITAL_ACT
   end for;
end CFG_IOIN_ID_VITAL;





---- CELL IOTRI_OD_EB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OD_EB is
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_E_EOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));




  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                E              :  in    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OD_EB :  entity is TRUE;
 end IOTRI_OD_EB;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OD_EB is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL DR_ipd  : STD_ULOGIC := 'X';
        SIGNAL DF_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
        SIGNAL OCLK_ipd : STD_ULOGIC := 'X';


 begin
         ---------------------
          --  INPUT PATH DELAYs
          ---------------------
          WireDelay : block
          begin
            VitalWireDelay (DR_ipd, DR, tipd_DR);
            VitalWireDelay (DF_ipd, DF, tipd_DF);
            VitalWireDelay (E_ipd,E, tipd_E);
            VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
            VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
          end block;



    --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (DR_ipd, DF_ipd,E_ipd,CLR_ipd,OCLK_ipd)

        -- timing check results
        VARIABLE Tviol_DR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_DF_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DF_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Pviol_OCLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_OCLK     : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_CLR      : STD_ULOGIC := '0';
        VARIABLE PInfo_CLR      : VitalPeriodDataType := VitalPeriodDataInit;

        -- functionality results
        VARIABLE Violation      : STD_ULOGIC := '0';
        VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE E_delayed    : STD_ULOGIC := 'X';
        VARIABLE DR_tmp    : STD_ULOGIC := 'X';
        VARIABLE DF_tmp    : STD_ULOGIC := 'X';

        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');

        ALIAS DOUT_zd : STD_LOGIC is Results(1);
        ALIAS EOUT_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
        VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

 begin

   ------------------------
   --  Timing Check Section
   ------------------------

   if(TimingChecksOn) then
        VitalSetupHoldCheck (
         Violation              => Tviol_DR_OCLK_posedge,
         TimingData             => Tmkr_DR_OCLK_posedge,
         TestSignal             => DR_ipd,
         TestSignalName         => "DR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DR_OCLK_posedge_posedge,
         SetupLow               => tsetup_DR_OCLK_negedge_posedge,
         HoldHigh               => thold_DR_OCLK_posedge_posedge,
         HoldLow                => thold_DR_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

         VitalSetupHoldCheck (
         Violation              => Tviol_DF_OCLK_posedge,
         TimingData             => Tmkr_DF_OCLK_posedge,
         TestSignal             => DF_ipd,
         TestSignalName         => "DF",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DF_OCLK_posedge_posedge,
         SetupLow               => tsetup_DF_OCLK_negedge_posedge,
         HoldHigh               => thold_DF_OCLK_posedge_posedge,
         HoldLow                => thold_DF_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);



      VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_OCLK_posedge,
         TimingData             => Tmkr_CLR_OCLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_OCLK_negedge_posedge,
         Removal               => thold_CLR_OCLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        VitalPeriodPulseCheck (
         Violation              => Pviol_OCLK,
         PeriodData             => PInfo_OCLK,
         TestSignal             => OCLK_ipd,
         TestSignalName         => "OCLK",
         TestDelay              => 0 ns,
         Period         => tperiod_OCLK_posedge,
         PulseWidthHigh => tpw_OCLK_posedge,
         PulseWidthLow => tpw_OCLK_negedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOTRI_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);



         VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period         => 0 ns,
         PulseWidthHigh => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOTRI_OD_EB",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        end if;




      --------------------------------
      --  Functionality Section
      -------------------------------

      Violation := Tviol_DR_OCLK_posedge or Tviol_DF_OCLK_posedge or Tviol_CLR_OCLK_posedge;

      VitalStateTable(
       Result => DR_tmp,
       PreviousDataIn => PrevData_QR,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DR_ipd ));
       DR_tmp := Violation XOR DR_tmp;

      VitalStateTable(
       Result => DF_tmp,
       PreviousDataIn => PrevData_QF,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DF_ipd ));
       DF_tmp := Violation XOR DF_tmp;

      DOUT_zd := VitalMUX2( DR_tmp, DF_tmp, OCLK_ipd );
      EOUT_zd := TO_X01( E_delayed );

      E_delayed  := E_ipd;



       ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
         OutSignal => DOUT,
         GlitchData => DOUT_GlitchData,
         OutSignalName => "DOUT",
         OutTemp => DOUT_zd,
         Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

       VitalPathDelay01 (
         OutSignal => EOUT,
         GlitchData => EOUT_GlitchData,
         OutSignalName => "EOUT",
         OutTemp => EOUT_zd,
         Paths => (0 => (E_ipd'last_event, tpd_E_EOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_IOTRI_OD_EB_VITAL of IOTRI_OD_EB is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OD_EB_VITAL;




---- CELL IOTRI_OD_ERC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOTRI_OD_ERC is
    generic(
                TimingChecksOn: Boolean := True;
                InstancePath: STRING := "*";
                Xon: Boolean := False;
                MsgOn: Boolean := True;
                tpd_CLR_DOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_DOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_CLR_EOUT      :  VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_OCLK_EOUT     :  VitalDelayType01 := (0.100 ns, 0.100 ns);

                tsetup_E_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_E_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DR_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;

                tsetup_DF_OCLK_posedge_posedge :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_posedge_posedge   :   VitalDelayType := 0.000 ns;
                tsetup_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                thold_DF_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;


                thold_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                trecovery_CLR_OCLK_negedge_posedge   :   VitalDelayType := 0.000 ns;
                tperiod_OCLK_posedge    :  VitalDelayType := 0.000 ns;
                tpw_OCLK_posedge :  VitalDelayType := 0.000 ns;
                tpw_OCLK_negedge  :  VitalDelayType := 0.000 ns;
                tpw_CLR_posedge :  VitalDelayType := 0.000 ns;
                tipd_DR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_DF        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_E        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_CLR        :   VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_OCLK            :    VitalDelayType01 := (0.000 ns, 0.000 ns));


  port(
                CLR             :   in    STD_ULOGIC;
                OCLK            :   in    STD_ULOGIC;
                DR             :  in    STD_ULOGIC;
                DF             :  in    STD_ULOGIC;
                E             :  in    STD_ULOGIC;
                DOUT               :  out    STD_ULOGIC;
                EOUT               :  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of IOTRI_OD_ERC :  entity is TRUE;
 end IOTRI_OD_ERC;







-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of IOTRI_OD_ERC is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL DR_ipd  : STD_ULOGIC := 'X';
        SIGNAL DF_ipd  : STD_ULOGIC := 'X';
        SIGNAL E_ipd  : STD_ULOGIC := 'X';
        SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
        SIGNAL OCLK_ipd : STD_ULOGIC := 'X';

begin

             ---------------------
             --  INPUT PATH DELAYs
             ---------------------
             WireDelay : block
             begin
               VitalWireDelay (DR_ipd, DR, tipd_DR);
               VitalWireDelay (DF_ipd, DF, tipd_DF);
               VitalWireDelay (E_ipd, E, tipd_E);
               VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
               VitalWireDelay (OCLK_ipd,OCLK, tipd_OCLK);
             end block;
  

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (DR_ipd, DF_ipd,E_ipd,CLR_ipd, OCLK_ipd)

        -- timing check results
        VARIABLE Tviol_DR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Tviol_DF_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_DF_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;

        VARIABLE Tviol_E_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_E_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;



        VARIABLE Tviol_CLR_OCLK_posedge         : STD_ULOGIC := '0';
        VARIABLE Tmkr_CLR_OCLK_posedge          : VitalTimingDataType := VitalTimingDataInit;
        VARIABLE Pviol_OCLK     : STD_ULOGIC := '0';
        VARIABLE PInfo_OCLK     : VitalPeriodDataType := VitalPeriodDataInit;
        VARIABLE Pviol_CLR      : STD_ULOGIC := '0';
        VARIABLE PInfo_CLR      : VitalPeriodDataType := VitalPeriodDataInit;

        -- functionality results
        VARIABLE Violation      : STD_ULOGIC := '0';
        VARIABLE PrevData_QE  : STD_LOGIC_VECTOR(0 to 6);
        VARIABLE PrevData_QR  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE PrevData_QF  : STD_LOGIC_VECTOR(0 to 2);
        VARIABLE OCLK_delayed   : STD_ULOGIC := 'X';
        VARIABLE E_delayed    : STD_ULOGIC := 'X';
        VARIABLE DR_tmp    : STD_ULOGIC := 'X';
        VARIABLE DF_tmp    : STD_ULOGIC := 'X';
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');

        ALIAS DOUT_zd : STD_LOGIC is Results(1);
        ALIAS EOUT_zd : STD_LOGIC is Results(2);

        -- output glitch detection variables
        VARIABLE DOUT_GlitchData  : VitalGlitchDataType;
        VARIABLE EOUT_GlitchData  : VitalGlitchDataType;

   begin

 
   ------------------------
   --  Timing Check Section
   ------------------------

   if(TimingChecksOn) then
        VitalSetupHoldCheck (
         Violation              => Tviol_DR_OCLK_posedge,
         TimingData             => Tmkr_DR_OCLK_posedge,
         TestSignal             => DR_ipd,
         TestSignalName         => "DR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DR_OCLK_posedge_posedge,
         SetupLow               => tsetup_DR_OCLK_negedge_posedge,
         HoldHigh               => thold_DR_OCLK_posedge_posedge,
         HoldLow                => thold_DR_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


         VitalSetupHoldCheck (
         Violation              => Tviol_DF_OCLK_posedge,
         TimingData             => Tmkr_DF_OCLK_posedge,
         TestSignal             => DF_ipd,
         TestSignalName         => "DF",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_DF_OCLK_posedge_posedge,
         SetupLow               => tsetup_DF_OCLK_negedge_posedge,
         HoldHigh               => thold_DF_OCLK_posedge_posedge,
         HoldLow                => thold_DF_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

        VitalSetupHoldCheck (
         Violation              => Tviol_E_OCLK_posedge,
         TimingData             => Tmkr_E_OCLK_posedge,
         TestSignal             => E_ipd,
         TestSignalName         => "E",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_E_OCLK_posedge_posedge,
         SetupLow               => tsetup_E_OCLK_negedge_posedge,
         HoldHigh               => thold_E_OCLK_posedge_posedge,
         HoldLow                => thold_E_OCLK_negedge_posedge,
         CheckEnabled           =>
            TO_X01((NOT CLR_ipd)) /= '0',
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);


        VitalRecoveryRemovalCheck (
         Violation              => Tviol_CLR_OCLK_posedge,
         TimingData             => Tmkr_CLR_OCLK_posedge,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         RefSignal              => OCLK_ipd,
         RefSignalName          => "OCLK",
         RefDelay               => 0 ns,
         Recovery              => trecovery_CLR_OCLK_negedge_posedge,
         Removal               => thold_CLR_OCLK_negedge_posedge,

         ActiveLow              => FALSE,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/IOTRI_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        VitalPeriodPulseCheck (
         Violation              => Pviol_OCLK,
         PeriodData             => PInfo_OCLK,
         TestSignal             => OCLK_ipd,
         TestSignalName         => "OCLK",
         TestDelay              => 0 ns,
         Period         => tperiod_OCLK_posedge,
         PulseWidthHigh => tpw_OCLK_posedge,
         PulseWidthLow => tpw_OCLK_negedge,
         CheckEnabled           =>
                TO_X01((( NOT CLR_ipd) ) ) /= '0',
         HeaderMsg              => InstancePath & "/IOTRI_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);


        VitalPeriodPulseCheck (
         Violation              => Pviol_CLR,
         PeriodData             => PInfo_CLR,
         TestSignal             => CLR_ipd,
         TestSignalName         => "CLR",
         TestDelay              => 0 ns,
         Period         => 0 ns,
         PulseWidthHigh => tpw_CLR_posedge,
         PulseWidthLow          => 0 ns,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/IOTRI_OD_ERC",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity            => WARNING);

        end if;

      --------------------------------
      --  Functionality Section
      -------------------------------

      Violation := Tviol_DR_OCLK_posedge or Tviol_E_OCLK_posedge or Tviol_DF_OCLK_posedge or Tviol_CLR_OCLK_posedge;

      VitalStateTable(
       Result => DR_tmp,
       PreviousDataIn => PrevData_QR,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DR_ipd ));
       DR_tmp := Violation XOR DR_tmp;

      VitalStateTable(
       Result => DF_tmp,
       PreviousDataIn => PrevData_QF,
       StateTable => DFN1C1_Q_tab,
       DataIn => ( CLR_ipd, OCLK_ipd, DF_ipd ));
       DF_tmp := Violation XOR DF_tmp;

      DOUT_zd := VitalMUX2( DR_tmp, DF_tmp, OCLK_ipd );

       VitalStateTable(
       Result => EOUT_zd,
       PreviousDataIn => PrevData_QE,
       StateTable => DFEG_Q_tab,
       DataIn => (
             (NOT CLR_ipd), OCLK_delayed, EOUT_zd, E_delayed,  '0', '1', OCLK_ipd));
       EOUT_zd := Violation XOR EOUT_zd;

      E_delayed  := E_ipd;
      OCLK_delayed :=OCLK_ipd;


      ----------------------
        --  Path Delay Section
        ----------------------
        VitalPathDelay01 (
         OutSignal => DOUT,
         GlitchData => DOUT_GlitchData,
         OutSignalName => "DOUT",
         OutTemp => DOUT_zd,
         Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_DOUT, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_DOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

       VitalPathDelay01 (
         OutSignal => EOUT,
         GlitchData => EOUT_GlitchData,
         OutSignalName => "EOUT",
         OutTemp => EOUT_zd,
         Paths => (0 => (OCLK_ipd'last_event, tpd_OCLK_EOUT, true),
                   1=> (CLR_ipd'last_event, tpd_CLR_EOUT, true)),
         Mode => OnDetect,
         Xon => Xon,
         MsgOn => MsgOn,
         MsgSeverity => WARNING);

   end process;

end VITAL_ACT;

configuration CFG_IOTRI_OD_ERC_VITAL of IOTRI_OD_ERC is
   for VITAL_ACT
   end for;
end CFG_IOTRI_OD_ERC_VITAL;



----- CELL RAM4K9 -----
library IEEE;
library STD;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_timing.all;
use IEEE.VITAL_primitives.all;


use std.textio.all;
use ieee.std_logic_textio.all;

 entity RAM4K9 is
   generic (
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;
      MEMORYFILE       : String  := "";
      WARNING_MSGS_ON  : Boolean := True;
           
      tipd_ADDRA11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRA0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB9      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB1      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ADDRB0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA8       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA7       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA6       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA5       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA4       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA3       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA2       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINA0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB8       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB7       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB6       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB5       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB4       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB3       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB2       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_DINB0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHA1     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHA0     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHB1     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WIDTHB0     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PIPEA       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PIPEB       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WMODEA      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WMODEB      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_BLKA        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_BLKB        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WENA        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WENB        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLKA        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLKB        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RESET       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLKA_DOUTA8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKA_DOUTA0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB8  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB7  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB6  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB5  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB4  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB3  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB2  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB1  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_CLKB_DOUTB0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA8 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA7 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA6 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA5 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA4 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA3 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA2 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA1 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTA0 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB8 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB7 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB6 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB5 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB4 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB3 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB2 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB1 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_DOUTB0 : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_DINA8_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA8_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA7_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA7_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA6_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA6_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA5_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA5_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA4_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA4_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA3_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA3_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA2_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA2_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA1_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA1_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA0_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINA0_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB8_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB8_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB7_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB7_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB6_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB6_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB5_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB5_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB4_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB4_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB3_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB3_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB2_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB2_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB1_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB1_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB0_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_DINB0_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_DINA8_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA8_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA7_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA7_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA6_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA6_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA5_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA5_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA4_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA4_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA3_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA3_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA2_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA2_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA1_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA1_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA0_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINA0_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB8_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB8_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB7_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB7_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB6_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB6_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB5_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB5_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB4_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB4_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB3_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB3_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB2_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB2_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB1_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB1_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB0_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_DINB0_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_ADDRA11_CLKA_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRA11_CLKA_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRA10_CLKA_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRA10_CLKA_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRA9_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA9_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA8_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA8_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA7_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA7_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA6_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA6_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA5_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA5_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA4_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA4_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA3_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA3_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA2_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA2_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA1_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA1_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA0_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRA0_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRA11_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRA11_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRA10_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRA10_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRA9_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA9_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA8_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA8_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA7_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA7_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA6_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA6_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA5_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA5_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA4_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA4_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA3_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA3_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA2_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA2_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA1_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA1_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA0_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRA0_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_ADDRB11_CLKB_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRB11_CLKB_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRB10_CLKB_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRB10_CLKB_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_ADDRB9_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB9_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB8_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB8_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB7_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB7_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB6_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB6_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB5_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB5_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB4_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB4_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB3_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB3_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB2_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB2_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB1_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB1_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB0_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_ADDRB0_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRB11_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRB11_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRB10_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRB10_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_ADDRB9_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB9_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB8_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB8_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB7_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB7_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB6_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB6_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB5_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB5_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB4_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB4_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB3_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB3_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB2_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB2_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB1_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB1_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB0_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_ADDRB0_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WENA_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WENA_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_BLKA_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_BLKA_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WMODEA_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WMODEA_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_PIPEA_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_PIPEA_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WENA_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WENA_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_BLKA_CLKA_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_BLKA_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WMODEA_CLKA_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WMODEA_CLKA_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_PIPEA_CLKA_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_PIPEA_CLKA_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WENB_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WENB_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_BLKB_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_BLKB_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WMODEB_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WMODEB_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_PIPEB_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_PIPEB_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB1_CLKB_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB1_CLKB_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_WIDTHB1_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHB1_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB0_CLKB_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WIDTHB0_CLKB_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_WIDTHB0_CLKB_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHB0_CLKB_posedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_WIDTHA1_CLKA_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WIDTHA1_CLKA_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_WIDTHA1_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHA1_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WIDTHA0_CLKA_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WIDTHA0_CLKA_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_WIDTHA0_CLKA_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WIDTHA0_CLKA_posedge_posedge  : VitalDelayType := 0.000 ns;

      thold_WENB_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WENB_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_BLKB_CLKB_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_BLKB_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WMODEB_CLKB_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WMODEB_CLKB_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_PIPEB_CLKB_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_PIPEB_CLKB_posedge_posedge    : VitalDelayType := 0.000 ns;
      
      tpw_CLKA_posedge                     : VitalDelayType := 0.000 ns;
      tpw_CLKA_negedge                     : VitalDelayType := 0.000 ns;
      tpw_CLKB_posedge                     : VitalDelayType := 0.000 ns;
      tpw_CLKB_negedge                     : VitalDelayType := 0.000 ns;
      trecovery_RESET_CLKA_posedge_posedge : VitalDelayType := 0.000 ns;
      trecovery_RESET_CLKB_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_RESET_CLKA_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RESET_CLKB_posedge_posedge     : VitalDelayType := 0.000 ns;
      tpw_RESET_negedge                    : VitalDelayType := 0.000 ns
     );

   port (
      ADDRA11       : IN STD_ULOGIC ;
      ADDRA10       : IN STD_ULOGIC ;
      ADDRA9        : IN STD_ULOGIC ;
      ADDRA8        : IN STD_ULOGIC ;
      ADDRA7        : IN STD_ULOGIC ;
      ADDRA6        : IN STD_ULOGIC ;
      ADDRA5        : IN STD_ULOGIC ;
      ADDRA4        : IN STD_ULOGIC ;
      ADDRA3        : IN STD_ULOGIC ;
      ADDRA2        : IN STD_ULOGIC ;
      ADDRA1        : IN STD_ULOGIC ;
      ADDRA0        : IN STD_ULOGIC ;
      ADDRB11       : IN STD_ULOGIC ;
      ADDRB10       : IN STD_ULOGIC ;
      ADDRB9        : IN STD_ULOGIC ;
      ADDRB8        : IN STD_ULOGIC ;
      ADDRB7        : IN STD_ULOGIC ;
      ADDRB6        : IN STD_ULOGIC ;
      ADDRB5        : IN STD_ULOGIC ;
      ADDRB4        : IN STD_ULOGIC ;
      ADDRB3        : IN STD_ULOGIC ;
      ADDRB2        : IN STD_ULOGIC ;
      ADDRB1        : IN STD_ULOGIC ;
      ADDRB0        : IN STD_ULOGIC ;
      DINA8         : IN STD_ULOGIC ;
      DINA7         : IN STD_ULOGIC ;
      DINA6         : IN STD_ULOGIC ;
      DINA5         : IN STD_ULOGIC ;
      DINA4         : IN STD_ULOGIC ;
      DINA3         : IN STD_ULOGIC ;
      DINA2         : IN STD_ULOGIC ;
      DINA1         : IN STD_ULOGIC ;
      DINA0         : IN STD_ULOGIC ; 
      DINB8         : IN STD_ULOGIC ;
      DINB7         : IN STD_ULOGIC ;
      DINB6         : IN STD_ULOGIC ;
      DINB5         : IN STD_ULOGIC ;
      DINB4         : IN STD_ULOGIC ;
      DINB3         : IN STD_ULOGIC ;
      DINB2         : IN STD_ULOGIC ;
      DINB1         : IN STD_ULOGIC ;
      DINB0         : IN STD_ULOGIC ;
      WIDTHA1       : IN STD_ULOGIC ;
      WIDTHA0       : IN STD_ULOGIC ;
      WIDTHB1       : IN STD_ULOGIC ;
      WIDTHB0       : IN STD_ULOGIC ;
      PIPEA         : IN STD_ULOGIC ;
      PIPEB         : IN STD_ULOGIC ;
      WMODEA        : IN STD_ULOGIC ;
      WMODEB        : IN STD_ULOGIC ;
      BLKA          : IN STD_ULOGIC ;
      BLKB          : IN STD_ULOGIC ;
      WENA          : IN STD_ULOGIC ;
      WENB          : IN STD_ULOGIC ;
      CLKA          : IN STD_ULOGIC ;
      CLKB          : IN STD_ULOGIC ;
      RESET         : IN STD_ULOGIC ;
      DOUTA8        : OUT STD_ULOGIC ;
      DOUTA7        : OUT STD_ULOGIC ;
      DOUTA6        : OUT STD_ULOGIC ;
      DOUTA5        : OUT STD_ULOGIC ;
      DOUTA4        : OUT STD_ULOGIC ;
      DOUTA3        : OUT STD_ULOGIC ;
      DOUTA2        : OUT STD_ULOGIC ;
      DOUTA1        : OUT STD_ULOGIC ;
      DOUTA0        : OUT STD_ULOGIC ;
      DOUTB8        : OUT STD_ULOGIC ;
      DOUTB7        : OUT STD_ULOGIC ;
      DOUTB6        : OUT STD_ULOGIC ;
      DOUTB5        : OUT STD_ULOGIC ;
      DOUTB4        : OUT STD_ULOGIC ;
      DOUTB3        : OUT STD_ULOGIC ;
      DOUTB2        : OUT STD_ULOGIC ;
      DOUTB1        : OUT STD_ULOGIC ;
      DOUTB0        : OUT STD_ULOGIC
     );
     
   attribute VITAL_LEVEL0 of RAM4K9 : entity is TRUE;

end RAM4K9;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4K9 is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;
  
  signal ADDRA11_ipd : std_ulogic := 'X';
  signal ADDRA10_ipd : std_ulogic := 'X';
  signal ADDRA9_ipd  : std_ulogic := 'X'; 
  signal ADDRA8_ipd  : std_ulogic := 'X';
  signal ADDRA7_ipd  : std_ulogic := 'X';
  signal ADDRA6_ipd  : std_ulogic := 'X'; 
  signal ADDRA5_ipd  : std_ulogic := 'X';
  signal ADDRA4_ipd  : std_ulogic := 'X';
  signal ADDRA3_ipd  : std_ulogic := 'X'; 
  signal ADDRA2_ipd  : std_ulogic := 'X';
  signal ADDRA1_ipd  : std_ulogic := 'X';
  signal ADDRA0_ipd  : std_ulogic := 'X'; 
  signal ADDRB11_ipd : std_ulogic := 'X';
  signal ADDRB10_ipd : std_ulogic := 'X';
  signal ADDRB9_ipd  : std_ulogic := 'X'; 
  signal ADDRB8_ipd  : std_ulogic := 'X';
  signal ADDRB7_ipd  : std_ulogic := 'X';
  signal ADDRB6_ipd  : std_ulogic := 'X'; 
  signal ADDRB5_ipd  : std_ulogic := 'X';
  signal ADDRB4_ipd  : std_ulogic := 'X';
  signal ADDRB3_ipd  : std_ulogic := 'X'; 
  signal ADDRB2_ipd  : std_ulogic := 'X';
  signal ADDRB1_ipd  : std_ulogic := 'X';
  signal ADDRB0_ipd  : std_ulogic := 'X'; 
  signal DINA8_ipd   : std_ulogic := 'X';
  signal DINA7_ipd   : std_ulogic := 'X';
  signal DINA6_ipd   : std_ulogic := 'X'; 
  signal DINA5_ipd   : std_ulogic := 'X';
  signal DINA4_ipd   : std_ulogic := 'X';
  signal DINA3_ipd   : std_ulogic := 'X'; 
  signal DINA2_ipd   : std_ulogic := 'X';
  signal DINA1_ipd   : std_ulogic := 'X';
  signal DINA0_ipd   : std_ulogic := 'X'; 
  signal DINB8_ipd   : std_ulogic := 'X';
  signal DINB7_ipd   : std_ulogic := 'X';
  signal DINB6_ipd   : std_ulogic := 'X'; 
  signal DINB5_ipd   : std_ulogic := 'X';
  signal DINB4_ipd   : std_ulogic := 'X';
  signal DINB3_ipd   : std_ulogic := 'X'; 
  signal DINB2_ipd   : std_ulogic := 'X';
  signal DINB1_ipd   : std_ulogic := 'X';
  signal DINB0_ipd   : std_ulogic := 'X'; 
  signal WIDTHA1_ipd : std_ulogic := 'X';
  signal WIDTHA0_ipd : std_ulogic := 'X'; 
  signal PIPEA_ipd   : std_ulogic := 'X';
  signal WMODEA_ipd  : std_ulogic := 'X';
  signal BLKA_ipd    : std_ulogic := 'X'; 
  signal WENA_ipd    : std_ulogic := 'X';
  signal CLKA_ipd    : std_ulogic := 'X';
  signal RESET_ipd   : std_ulogic := 'X'; 
  signal WIDTHB1_ipd : std_ulogic := 'X';
  signal WIDTHB0_ipd : std_ulogic := 'X'; 
  signal PIPEB_ipd   : std_ulogic := 'X';
  signal WMODEB_ipd  : std_ulogic := 'X';
  signal BLKB_ipd    : std_ulogic := 'X'; 
  signal WENB_ipd    : std_ulogic := 'X';
  signal CLKB_ipd    : std_ulogic := 'X';
  
  signal INIT_MEM    : std_logic  := '0';

  type MEMORY_512_9 is array ( 0 to 511, 8 downto 0 ) of std_ulogic; -- memory array with pre-load capability

  constant TC2CWRH   : time       := 1.013 ns;
  constant TC2CRWH   : time       := 0.883 ns;
  constant TC2CWWL   : time       := 0.3 ns;

  -- 
  -- function to check if write and read operations are accessing the same memory location
  -- 

  function same_addr(
    waddr, raddr : integer;
    ww, rw       : integer ) return boolean is
    variable result           : boolean;
    variable wr_addr, rd_addr : integer;
  begin
    result := false;

    if ( ww > rw ) then
      rd_addr := ( raddr / (2 ** (ww-rw)) );
      wr_addr := waddr;
    elsif ( rw > ww ) then
      rd_addr := raddr;
      wr_addr := ( waddr / (2 ** (rw-ww)) );
    else
      rd_addr := raddr;
      wr_addr := waddr;
    end if;

    if ( wr_addr = rd_addr ) then
      result := true;
    end if;

    return result;
  end function same_addr;

  -- 
  -- function to drive read data bus to "x" depending on width configuration
  -- 

  function drive_data_x(
    waddr, raddr : integer;
    ww, rw       : integer;
    rd_data      : std_logic_vector (8 downto 0) ) return std_logic_vector is

    variable data_x : std_logic_vector (8 downto 0);
    variable index  : integer;

  begin
    data_x := rd_data;

    case (rw) is
      when 0 =>
            data_x (0) := 'X';
      when 1 =>
            if ( ww = 0 ) then
              data_x ( waddr mod 2 ) := 'X';
            else
              data_x ( 1 downto 0 ) := ( others => 'X' );
            end if;
      when 2 =>
            if ( ww = 0 ) then
              data_x ( waddr mod 4 ) := 'X';
            elsif ( ww = 1 ) then
              index := ( waddr mod 2 ) * 2;
              for i in index to index+1 loop
                data_x ( i ) := 'X';
              end loop;
            else
              data_x ( 3 downto 0 ) := ( others => 'X' );
            end if;
      when 3 =>
            if ( ww = 0 ) then
              data_x ( ( waddr mod 8 ) ) := 'X';
            elsif ( ww = 1 ) then
              index := ( waddr mod 4 ) * 2;
              for i in index to index+1 loop
                data_x ( i ) := 'X';
              end loop;
            elsif ( ww = 2 ) then
              index := ( waddr mod 2 ) * 4;
              for i in index to index+3 loop
                data_x ( i ) := 'X';
              end loop;
            else
              data_x ( 8 downto 0 ) := ( others => 'X' );
            end if;
      when others =>
            assert false
              report ": Invalid READ WIDTH, Legal Width: 0,1,2,3"
              severity warning;

     end case;

    return data_x;

  end function drive_data_x;


  begin  --  VITAL_ACT

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WireDelay: block

  begin  --  block WireDelay
    VitalWireDelay ( ADDRA11_ipd, ADDRA11, VitalExtendToFillDelay(tipd_ADDRA11) );
    VitalWireDelay ( ADDRA10_ipd, ADDRA10, VitalExtendToFillDelay(tipd_ADDRA10) );
    VitalWireDelay ( ADDRA9_ipd,  ADDRA9,  VitalExtendToFillDelay(tipd_ADDRA9)  );
    VitalWireDelay ( ADDRA8_ipd,  ADDRA8,  VitalExtendToFillDelay(tipd_ADDRA8)  );
    VitalWireDelay ( ADDRA7_ipd,  ADDRA7,  VitalExtendToFillDelay(tipd_ADDRA7)  );
    VitalWireDelay ( ADDRA6_ipd,  ADDRA6,  VitalExtendToFillDelay(tipd_ADDRA6)  );
    VitalWireDelay ( ADDRA5_ipd,  ADDRA5,  VitalExtendToFillDelay(tipd_ADDRA5)  );
    VitalWireDelay ( ADDRA4_ipd,  ADDRA4,  VitalExtendToFillDelay(tipd_ADDRA4)  );
    VitalWireDelay ( ADDRA3_ipd,  ADDRA3,  VitalExtendToFillDelay(tipd_ADDRA3)  );
    VitalWireDelay ( ADDRA2_ipd,  ADDRA2,  VitalExtendToFillDelay(tipd_ADDRA2)  );
    VitalWireDelay ( ADDRA1_ipd,  ADDRA1,  VitalExtendToFillDelay(tipd_ADDRA1)  );
    VitalWireDelay ( ADDRA0_ipd,  ADDRA0,  VitalExtendToFillDelay(tipd_ADDRA0)  );
    VitalWireDelay ( ADDRB11_ipd, ADDRB11, VitalExtendToFillDelay(tipd_ADDRB11) );
    VitalWireDelay ( ADDRB10_ipd, ADDRB10, VitalExtendToFillDelay(tipd_ADDRB10) );
    VitalWireDelay ( ADDRB9_ipd,  ADDRB9,  VitalExtendToFillDelay(tipd_ADDRB9)  );
    VitalWireDelay ( ADDRB8_ipd,  ADDRB8,  VitalExtendToFillDelay(tipd_ADDRB8)  );
    VitalWireDelay ( ADDRB7_ipd,  ADDRB7,  VitalExtendToFillDelay(tipd_ADDRB7)  );
    VitalWireDelay ( ADDRB6_ipd,  ADDRB6,  VitalExtendToFillDelay(tipd_ADDRB6)  );
    VitalWireDelay ( ADDRB5_ipd,  ADDRB5,  VitalExtendToFillDelay(tipd_ADDRB5)  );
    VitalWireDelay ( ADDRB4_ipd,  ADDRB4,  VitalExtendToFillDelay(tipd_ADDRB4)  );
    VitalWireDelay ( ADDRB3_ipd,  ADDRB3,  VitalExtendToFillDelay(tipd_ADDRB3)  );
    VitalWireDelay ( ADDRB2_ipd,  ADDRB2,  VitalExtendToFillDelay(tipd_ADDRB2)  );
    VitalWireDelay ( ADDRB1_ipd,  ADDRB1,  VitalExtendToFillDelay(tipd_ADDRB1)  );
    VitalWireDelay ( ADDRB0_ipd,  ADDRB0,  VitalExtendToFillDelay(tipd_ADDRB0)  );
    VitalWireDelay ( DINA8_ipd,   DINA8,   VitalExtendToFillDelay(tipd_DINA8)   );
    VitalWireDelay ( DINA7_ipd,   DINA7,   VitalExtendToFillDelay(tipd_DINA7)   );
    VitalWireDelay ( DINA6_ipd,   DINA6,   VitalExtendToFillDelay(tipd_DINA6)   );
    VitalWireDelay ( DINA5_ipd,   DINA5,   VitalExtendToFillDelay(tipd_DINA5)   );
    VitalWireDelay ( DINA4_ipd,   DINA4,   VitalExtendToFillDelay(tipd_DINA4)   );
    VitalWireDelay ( DINA3_ipd,   DINA3,   VitalExtendToFillDelay(tipd_DINA3)   );
    VitalWireDelay ( DINA2_ipd,   DINA2,   VitalExtendToFillDelay(tipd_DINA2)   );
    VitalWireDelay ( DINA1_ipd,   DINA1,   VitalExtendToFillDelay(tipd_DINA1)   );
    VitalWireDelay ( DINA0_ipd,   DINA0,   VitalExtendToFillDelay(tipd_DINA0)   );
    VitalWireDelay ( DINB8_ipd,   DINB8,   VitalExtendToFillDelay(tipd_DINB8)   );
    VitalWireDelay ( DINB7_ipd,   DINB7,   VitalExtendToFillDelay(tipd_DINB7)   );
    VitalWireDelay ( DINB6_ipd,   DINB6,   VitalExtendToFillDelay(tipd_DINB6)   );
    VitalWireDelay ( DINB5_ipd,   DINB5,   VitalExtendToFillDelay(tipd_DINB5)   );
    VitalWireDelay ( DINB4_ipd,   DINB4,   VitalExtendToFillDelay(tipd_DINB4)   );
    VitalWireDelay ( DINB3_ipd,   DINB3,   VitalExtendToFillDelay(tipd_DINB3)   );
    VitalWireDelay ( DINB2_ipd,   DINB2,   VitalExtendToFillDelay(tipd_DINB2)   );
    VitalWireDelay ( DINB1_ipd,   DINB1,   VitalExtendToFillDelay(tipd_DINB1)   );
    VitalWireDelay ( DINB0_ipd,   DINB0,   VitalExtendToFillDelay(tipd_DINB0)   );
    VitalWireDelay ( WIDTHA1_ipd, WIDTHA1, VitalExtendToFillDelay(tipd_WIDTHA1) );
    VitalWireDelay ( WIDTHA0_ipd, WIDTHA0, VitalExtendToFillDelay(tipd_WIDTHA0) );
    VitalWireDelay ( PIPEA_ipd,   PIPEA,   VitalExtendToFillDelay(tipd_PIPEA)   );
    VitalWireDelay ( WMODEA_ipd,  WMODEA,  VitalExtendToFillDelay(tipd_WMODEA)  );
    VitalWireDelay ( BLKA_ipd,    BLKA,    VitalExtendToFillDelay(tipd_BLKA)    );
    VitalWireDelay ( WENA_ipd,    WENA,    VitalExtendToFillDelay(tipd_WENA)    );
    VitalWireDelay ( CLKA_ipd,    CLKA,    VitalExtendToFillDelay(tipd_CLKA)    );
    VitalWireDelay ( WIDTHB1_ipd, WIDTHB1, VitalExtendToFillDelay(tipd_WIDTHB1) );
    VitalWireDelay ( WIDTHB0_ipd, WIDTHB0, VitalExtendToFillDelay(tipd_WIDTHB0) );
    VitalWireDelay ( PIPEB_ipd,   PIPEB,   VitalExtendToFillDelay(tipd_PIPEB)   );
    VitalWireDelay ( WMODEB_ipd,  WMODEB,  VitalExtendToFillDelay(tipd_WMODEB)  );
    VitalWireDelay ( BLKB_ipd,    BLKB,    VitalExtendToFillDelay(tipd_BLKB)    );
    VitalWireDelay ( WENB_ipd,    WENB,    VitalExtendToFillDelay(tipd_WENB)    );
    VitalWireDelay ( CLKB_ipd,    CLKB,    VitalExtendToFillDelay(tipd_CLKB)    );
    VitalWireDelay ( RESET_ipd,   RESET,   VitalExtendToFillDelay(tipd_RESET)   );
   
  end block WireDelay;

  -- INITIALIZE MEMORY --

  process
  begin
    INIT_MEM <= '1';
    wait;
  end process;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (CLKA_ipd, WENA_ipd, PIPEA_ipd, WIDTHA1_ipd, WIDTHA0_ipd, 
                           BLKA_ipd, WMODEA_ipd, RESET_ipd,
                           CLKB_ipd, WENB_ipd, PIPEB_ipd, WIDTHB1_ipd, WIDTHB0_ipd,
                           BLKB_ipd, WMODEB_ipd,
                           ADDRA11_ipd, ADDRA10_ipd, ADDRA9_ipd, ADDRA8_ipd, 
                           ADDRA7_ipd, ADDRA6_ipd, ADDRA5_ipd, ADDRA4_ipd,
                           ADDRA3_ipd, ADDRA2_ipd, ADDRA1_ipd, ADDRA0_ipd, 
                           ADDRB11_ipd, ADDRB10_ipd, ADDRB9_ipd, ADDRB8_ipd,
                           ADDRB7_ipd, ADDRB6_ipd, ADDRB5_ipd, ADDRB4_ipd,
                           ADDRB3_ipd, ADDRB2_ipd, ADDRB1_ipd, ADDRB0_ipd,
                           DINA8_ipd, DINA7_ipd, DINA6_ipd, DINA5_ipd, DINA4_ipd,
                           DINA3_ipd, DINA2_ipd, DINA1_ipd, DINA0_ipd,
                           DINB8_ipd, DINB7_ipd, DINB6_ipd, DINB5_ipd, DINB4_ipd,
                           DINB3_ipd, DINB2_ipd, DINB1_ipd, DINB0_ipd, INIT_MEM
                          )


     -- some internal veriable declaration
     variable ADDRA  : integer := 0;
     variable ADDRB  : integer := 0;
     variable widthA : integer := 0;
     variable widthB : integer := 0;

     variable ADDRA_VALID : integer := 1;
     variable ADDRB_VALID : integer := 1;

     variable MEM_512_9 : MEMORY_512_9;

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);

     variable i              : integer := 0;
     file     memfile        : text;
     variable status         : file_open_status;
     variable msgs_checked   : Boolean := False;
 
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-4095, -4095, 0, 1, -4095, -4095, 0, 1, -4095);

     --  Read Timing Check Results
     variable Tviol_DINA8_CLKA_posedge : X01 := '0';
     variable TmDt_DINA8_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA7_CLKA_posedge : X01 := '0';
     variable TmDt_DINA7_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA6_CLKA_posedge : X01 := '0';
     variable TmDt_DINA6_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA5_CLKA_posedge : X01 := '0';
     variable TmDt_DINA5_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA4_CLKA_posedge : X01 := '0';
     variable TmDt_DINA4_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA3_CLKA_posedge : X01 := '0';
     variable TmDt_DINA3_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA2_CLKA_posedge : X01 := '0';
     variable TmDt_DINA2_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA1_CLKA_posedge : X01 := '0';
     variable TmDt_DINA1_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINA0_CLKA_posedge : X01 := '0';
     variable TmDt_DINA0_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB8_CLKB_posedge : X01 := '0';
     variable TmDt_DINB8_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB7_CLKB_posedge : X01 := '0';
     variable TmDt_DINB7_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB6_CLKB_posedge : X01 := '0';
     variable TmDt_DINB6_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB5_CLKB_posedge : X01 := '0';
     variable TmDt_DINB5_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB4_CLKB_posedge : X01 := '0';
     variable TmDt_DINB4_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB3_CLKB_posedge : X01 := '0';
     variable TmDt_DINB3_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB2_CLKB_posedge : X01 := '0';
     variable TmDt_DINB2_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB1_CLKB_posedge : X01 := '0';
     variable TmDt_DINB1_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DINB0_CLKB_posedge : X01 := '0';
     variable TmDt_DINB0_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;

     variable Tviol_ADDRA11_CLKA_posedge : X01 := '0';
     variable TmDt_ADDRA11_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA10_CLKA_posedge : X01 := '0';
     variable TmDt_ADDRA10_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA9_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA9_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA8_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA8_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA7_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA7_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA6_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA6_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA5_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA5_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA4_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA4_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA3_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA3_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA2_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA2_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA1_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA1_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRA0_CLKA_posedge  : X01 := '0';
     variable TmDt_ADDRA0_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
    
     variable Tviol_ADDRB11_CLKB_posedge : X01 := '0';
     variable TmDt_ADDRB11_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB10_CLKB_posedge : X01 := '0';
     variable TmDt_ADDRB10_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB9_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB9_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB8_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB8_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB7_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB7_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB6_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB6_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB5_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB5_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB4_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB4_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB3_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB3_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB2_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB2_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB1_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB1_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ADDRB0_CLKB_posedge  : X01 := '0';
     variable TmDt_ADDRB0_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
    
     variable Tviol_WIDTHA1_CLKA_posedge : X01 := '0';
     variable TmDt_WIDTHA1_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTHA0_CLKA_posedge : X01 := '0';
     variable TmDt_WIDTHA0_CLKA_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PIPEA_CLKA_posedge   : X01 := '0';
     variable TmDt_PIPEA_CLKA_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WMODEA_CLKA_posedge  : X01 := '0';
     variable TmDt_WMODEA_CLKA_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKA_CLKA_posedge    : X01 := '0';
     variable TmDt_BLKA_CLKA_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENA_CLKA_posedge    : X01 := '0';
     variable TmDt_WENA_CLKA_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTHB1_CLKB_posedge : X01 := '0';
     variable TmDt_WIDTHB1_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WIDTHB0_CLKB_posedge : X01 := '0';
     variable TmDt_WIDTHB0_CLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PIPEB_CLKB_posedge   : X01 := '0';
     variable TmDt_PIPEB_CLKB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WMODEB_CLKB_posedge  : X01 := '0';
     variable TmDt_WMODEB_CLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKB_CLKB_posedge    : X01 := '0';
     variable TmDt_BLKB_CLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WENB_CLKB_posedge    : X01 := '0';
     variable TmDt_WENB_CLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
 
     variable Pviol_CLKA                 : X01 := '0';
     variable PeriodData_CLKA            : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_CLKB                 : X01 := '0';
     variable PeriodData_CLKB            : VitalPeriodDataType := VitalPeriodDataInit;
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01 := '0';
     variable Tviol_RESET_CLKA_posedge   : X01 := '0';
     variable Tmkr_RESET_CLKA_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_CLKB_posedge   : X01 := '0';
     variable Tmkr_RESET_CLKB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLKA_CLKB_posedge    : X01 := '0';
     variable TmDt_CLKA_CLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_CLKB_CLKA_posedge    : X01 := '0';
     variable TmDt_CLKB_CLKA_posedge     : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable DOUTA8_zd : std_ulogic;
     variable DOUTA7_zd : std_ulogic;
     variable DOUTA6_zd : std_ulogic;
     variable DOUTA5_zd : std_ulogic;
     variable DOUTA4_zd : std_ulogic;
     variable DOUTA3_zd : std_ulogic;
     variable DOUTA2_zd : std_ulogic;
     variable DOUTA1_zd : std_ulogic;
     variable DOUTA0_zd : std_ulogic;
     variable DOUTB8_zd : std_ulogic; 
     variable DOUTB7_zd : std_ulogic;
     variable DOUTB6_zd : std_ulogic;
     variable DOUTB5_zd : std_ulogic;
     variable DOUTB4_zd : std_ulogic;
     variable DOUTB3_zd : std_ulogic;
     variable DOUTB2_zd : std_ulogic;
     variable DOUTB1_zd : std_ulogic;
     variable DOUTB0_zd : std_ulogic;

     variable DOUTA8_stg : std_ulogic;
     variable DOUTA7_stg : std_ulogic;
     variable DOUTA6_stg : std_ulogic;
     variable DOUTA5_stg : std_ulogic;
     variable DOUTA4_stg : std_ulogic;
     variable DOUTA3_stg : std_ulogic;
     variable DOUTA2_stg : std_ulogic;
     variable DOUTA1_stg : std_ulogic;
     variable DOUTA0_stg : std_ulogic;
     variable DOUTB8_stg : std_ulogic;
     variable DOUTB7_stg : std_ulogic;
     variable DOUTB6_stg : std_ulogic;
     variable DOUTB5_stg : std_ulogic;
     variable DOUTB4_stg : std_ulogic;
     variable DOUTB3_stg : std_ulogic;
     variable DOUTB2_stg : std_ulogic;
     variable DOUTB1_stg : std_ulogic;
     variable DOUTB0_stg : std_ulogic;

     -- Output Glitch Detection Support Variables

     variable DOUTA8_GlitchData : VitalGlitchDataType;
     variable DOUTA7_GlitchData : VitalGlitchDataType;
     variable DOUTA6_GlitchData : VitalGlitchDataType;
     variable DOUTA5_GlitchData : VitalGlitchDataType;
     variable DOUTA4_GlitchData : VitalGlitchDataType;
     variable DOUTA3_GlitchData : VitalGlitchDataType;
     variable DOUTA2_GlitchData : VitalGlitchDataType;
     variable DOUTA1_GlitchData : VitalGlitchDataType;
     variable DOUTA0_GlitchData : VitalGlitchDataType;
     variable DOUTB8_GlitchData : VitalGlitchDataType;
     variable DOUTB7_GlitchData : VitalGlitchDataType;
     variable DOUTB6_GlitchData : VitalGlitchDataType;
     variable DOUTB5_GlitchData : VitalGlitchDataType;
     variable DOUTB4_GlitchData : VitalGlitchDataType;
     variable DOUTB3_GlitchData : VitalGlitchDataType;
     variable DOUTB2_GlitchData : VitalGlitchDataType;
     variable DOUTB1_GlitchData : VitalGlitchDataType;
     variable DOUTB0_GlitchData : VitalGlitchDataType;

      -- last value variables
      
     variable CLKA_previous : std_ulogic := 'X';
     variable CLKB_previous : std_ulogic := 'X';

     variable WENA_delayed  : std_ulogic := 'X';
     variable WENB_delayed  : std_ulogic := 'X';
     variable PIPEA_delayed : std_ulogic := 'X';
     variable PIPEB_delayed : std_ulogic := 'X';
     variable RESET_delayed : std_ulogic := 'X';
     variable BLKB_delayed  : std_ulogic := 'X';
     variable BLKA_delayed  : std_ulogic := 'X';
 

     variable ADDRA11_delayed : std_ulogic := 'X';
     variable ADDRA10_delayed : std_ulogic := 'X';  
     variable ADDRA9_delayed  : std_ulogic := 'X';
     variable ADDRA8_delayed  : std_ulogic := 'X';
     variable ADDRA7_delayed  : std_ulogic := 'X';
     variable ADDRA6_delayed  : std_ulogic := 'X';
     variable ADDRA5_delayed  : std_ulogic := 'X';
     variable ADDRA4_delayed  : std_ulogic := 'X';
     variable ADDRA3_delayed  : std_ulogic := 'X';
     variable ADDRA2_delayed  : std_ulogic := 'X';
     variable ADDRA1_delayed  : std_ulogic := 'X';
     variable ADDRA0_delayed  : std_ulogic := 'X';

     variable ADDRB11_delayed : std_ulogic := 'X';  
     variable ADDRB10_delayed : std_ulogic := 'X';  
     variable ADDRB9_delayed  : std_ulogic := 'X';
     variable ADDRB8_delayed  : std_ulogic := 'X';
     variable ADDRB7_delayed  : std_ulogic := 'X';
     variable ADDRB6_delayed  : std_ulogic := 'X';
     variable ADDRB5_delayed  : std_ulogic := 'X';
     variable ADDRB4_delayed  : std_ulogic := 'X';
     variable ADDRB3_delayed  : std_ulogic := 'X';
     variable ADDRB2_delayed  : std_ulogic := 'X';
     variable ADDRB1_delayed  : std_ulogic := 'X';
     variable ADDRB0_delayed  : std_ulogic := 'X';

     variable DINA8_delayed   : std_ulogic := 'X';
     variable DINA7_delayed   : std_ulogic := 'X';
     variable DINA6_delayed   : std_ulogic := 'X';
     variable DINA5_delayed   : std_ulogic := 'X';
     variable DINA4_delayed   : std_ulogic := 'X';
     variable DINA3_delayed   : std_ulogic := 'X';
     variable DINA2_delayed   : std_ulogic := 'X';
     variable DINA1_delayed   : std_ulogic := 'X';
     variable DINA0_delayed   : std_ulogic := 'X';

     variable DINB8_delayed   : std_ulogic := 'X';
     variable DINB7_delayed   : std_ulogic := 'X';
     variable DINB6_delayed   : std_ulogic := 'X';
     variable DINB5_delayed   : std_ulogic := 'X';
     variable DINB4_delayed   : std_ulogic := 'X';
     variable DINB3_delayed   : std_ulogic := 'X';
     variable DINB2_delayed   : std_ulogic := 'X';
     variable DINB1_delayed   : std_ulogic := 'X';
     variable DINB0_delayed   : std_ulogic := 'X';

     -- simultaneous write and read logic detection

     variable WENA_lat        : std_logic;
     variable WENB_lat        : std_logic;
     variable WDA_INT         : integer := 0;
     variable WDB_INT         : integer := 0;
     variable CLKA_wr_re      : Time;
     variable CLKA_wr_fe      : Time;
     variable CLKA_rd_re      : Time;
     variable CLKB_wr_re      : Time;
     variable CLKB_wr_fe      : Time;
     variable CLKB_rd_re      : Time;
     variable DOUTA_array     : std_logic_vector ( 8 downto 0 );
     variable DOUTB_array     : std_logic_vector ( 8 downto 0 );
     variable DINA_array      : std_logic_vector ( 8 downto 0 );
     variable DINB_array      : std_logic_vector ( 8 downto 0 );
 
     variable DINA8_bypass    : std_logic;
     variable DINA7_bypass    : std_logic;
     variable DINA6_bypass    : std_logic;
     variable DINA5_bypass    : std_logic;
     variable DINA4_bypass    : std_logic;
     variable DINA3_bypass    : std_logic;
     variable DINA2_bypass    : std_logic;
     variable DINA1_bypass    : std_logic;
     variable DINA0_bypass    : std_logic;

     variable DINB8_bypass    : std_logic;
     variable DINB7_bypass    : std_logic;
     variable DINB6_bypass    : std_logic;
     variable DINB5_bypass    : std_logic;
     variable DINB4_bypass    : std_logic;
     variable DINB3_bypass    : std_logic;
     variable DINB2_bypass    : std_logic;
     variable DINB1_bypass    : std_logic;
     variable DINB0_bypass    : std_logic;

begin -- process VITALBehavior

  if ( msgs_checked = False ) then
    msgs_checked := True;
    if ( WARNING_MSGS_ON = False ) then
      report "RAM4K9 warnings disabled. Set WARNING_MSGS_ON => True to enable."
      severity note;
    end if;
  end if;
  
  
  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------
  
  if ( INIT_MEM'event and INIT_MEM = '1' ) then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while (( i <= 511 ) and ( not endfile(memfile))) loop
        readline(memfile, inline);
        read(inline, indata);
        resdata := indata;
        MEM_512_9(i,8) := resdata(8);
        MEM_512_9(i,7) := resdata(7);
        MEM_512_9(i,6) := resdata(6);
        MEM_512_9(i,5) := resdata(5);
        MEM_512_9(i,4) := resdata(4);
        MEM_512_9(i,3) := resdata(3);
        MEM_512_9(i,2) := resdata(2);
        MEM_512_9(i,1) := resdata(1);
        MEM_512_9(i,0) := resdata(0);
        i := i + 1;
      end loop;
    else
      if ( WARNING_MSGS_ON ) then
        assert ( MEMORYFILE'length = 0 )
          report "Failed to open memory initialization in read mode"
          severity note;
      end if;
    end if;
    file_close(memfile);
  end if;


  if (TimingChecksOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery/ removal check for CLKA to RESET signal ;
     VitalRecoveryRemovalCheck   (
         Violation              => Tviol_RESET_CLKA_posedge,
         TimingData             => Tmkr_RESET_CLKA_posedge,
         TestSignal             => RESET_ipd,
         TestSignalName         => "RESET",
         TestDelay              => 0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0 ns,
         Recovery               => trecovery_RESET_CLKA_posedge_posedge,
         Removal                => thold_RESET_CLKA_posedge_posedge,
         ActiveLow              => TRUE,
         CheckEnabled           => (TO_X01(BLKA_ipd) = '0'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

    -- recovery/ removal check for CLKB to RESET signal ;
     VitalRecoveryRemovalCheck   (
         Violation              => Tviol_RESET_CLKB_posedge,
         TimingData             => Tmkr_RESET_CLKB_posedge,
         TestSignal             => RESET_ipd,
         TestSignalName         => "RESET",
         TestDelay              => 0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0 ns,
         Recovery               => trecovery_RESET_CLKB_posedge_posedge,
         Removal                => thold_RESET_CLKB_posedge_posedge,
         ActiveLow              => TRUE,
         CheckEnabled           => (TO_X01(BLKB_ipd) = '0'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

    -- setup / hold WENA to CLKA
     VitalSetupHoldCheck (
         Violation              => Tviol_WENA_CLKA_posedge,
         TimingData             => TmDt_WENA_CLKA_posedge,
         TestSignal             => WENA_ipd,
         TestSignalName         => "WENA",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WENA_CLKA_posedge_posedge,
         SetupLow               => tsetup_WENA_CLKA_negedge_posedge,
         HoldHigh               => thold_WENA_CLKA_posedge_posedge,
         HoldLow                => thold_WENA_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_PIPEA_CLKA_posedge,
         TimingData             => TmDt_PIPEA_CLKA_posedge,
         TestSignal             => PIPEA_ipd, 
         TestSignalName         => "PIPEA",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_PIPEA_CLKA_posedge_posedge,
         SetupLow               => tsetup_PIPEA_CLKA_negedge_posedge,
         HoldHigh               => thold_PIPEA_CLKA_posedge_posedge,
         HoldLow                => thold_PIPEA_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_BLKA_CLKA_posedge,
         TimingData             => TmDt_BLKA_CLKA_posedge,
         TestSignal             => BLKA_ipd, 
         TestSignalName         => "BLKA",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_BLKA_CLKA_posedge_posedge,
         SetupLow               => tsetup_BLKA_CLKA_negedge_posedge,
         HoldHigh               => thold_BLKA_CLKA_posedge_posedge,
         HoldLow                => thold_BLKA_CLKA_negedge_posedge,
         CheckEnabled           => (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WENB_CLKB_posedge,
         TimingData             => TmDt_WENB_CLKB_posedge,
         TestSignal             => WENB_ipd, 
         TestSignalName         => "WENB",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WENB_CLKB_posedge_posedge,
         SetupLow               => tsetup_WENB_CLKB_negedge_posedge,
         HoldHigh               => thold_WENB_CLKB_posedge_posedge,
         HoldLow                => thold_WENB_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_PIPEB_CLKB_posedge,
         TimingData             => TmDt_PIPEB_CLKB_posedge,
         TestSignal             => PIPEB_ipd, 
         TestSignalName         => "PIPEB",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_PIPEB_CLKB_posedge_posedge,
         SetupLow               => tsetup_PIPEB_CLKB_negedge_posedge,
         HoldHigh               => thold_PIPEB_CLKB_posedge_posedge,
         HoldLow                => thold_PIPEB_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_BLKB_CLKB_posedge,
         TimingData             => TmDt_BLKB_CLKB_posedge,
         TestSignal             => BLKB_ipd, 
         TestSignalName         => "BLKB",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_BLKB_CLKB_posedge_posedge,
         SetupLow               => tsetup_BLKB_CLKB_negedge_posedge,
         HoldHigh               => thold_BLKB_CLKB_posedge_posedge,
         HoldLow                => thold_BLKB_CLKB_negedge_posedge,
         CheckEnabled           => (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WIDTHB1_CLKB_posedge,
         TimingData             => TmDt_WIDTHB1_CLKB_posedge,
         TestSignal             => WIDTHB1_ipd, 
         TestSignalName         => "WIDTHB1",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WIDTHB1_CLKB_posedge_posedge,
         SetupLow               => tsetup_WIDTHB1_CLKB_negedge_posedge,
         HoldHigh               => thold_WIDTHB1_CLKB_posedge_posedge,
         HoldLow                => thold_WIDTHB1_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WIDTHB0_CLKB_posedge,
         TimingData             => TmDt_WIDTHB0_CLKB_posedge,
         TestSignal             => WIDTHB0_ipd, 
         TestSignalName         => "WIDTHB0",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WIDTHB0_CLKB_posedge_posedge,
         SetupLow               => tsetup_WIDTHB0_CLKB_negedge_posedge,
         HoldHigh               => thold_WIDTHB0_CLKB_posedge_posedge,
         HoldLow                => thold_WIDTHB0_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WMODEB_CLKB_posedge,
         TimingData             => TmDt_WMODEB_CLKB_posedge,
         TestSignal             => WMODEB_ipd, 
         TestSignalName         => "WMODEB",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WMODEB_CLKB_posedge_posedge,
         SetupLow               => tsetup_WMODEB_CLKB_negedge_posedge,
         HoldHigh               => thold_WMODEB_CLKB_posedge_posedge,
         HoldLow                => thold_WMODEB_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WIDTHA1_CLKA_posedge,
         TimingData             => TmDt_WIDTHA1_CLKA_posedge,
         TestSignal             => WIDTHA1_ipd, 
         TestSignalName         => "WIDTHA1",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WIDTHA1_CLKA_posedge_posedge,
         SetupLow               => tsetup_WIDTHA1_CLKA_negedge_posedge,
         HoldHigh               => thold_WIDTHA1_CLKA_posedge_posedge,
         HoldLow                => thold_WIDTHA1_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WIDTHA0_CLKA_posedge,
         TimingData             => TmDt_WIDTHA0_CLKA_posedge,
         TestSignal             => WIDTHA0_ipd, 
         TestSignalName         => "WIDTHA0",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WIDTHA0_CLKA_posedge_posedge,
         SetupLow               => tsetup_WIDTHA0_CLKA_negedge_posedge,
         HoldHigh               => thold_WIDTHA0_CLKA_posedge_posedge,
         HoldLow                => thold_WIDTHA0_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_WMODEA_CLKA_posedge,
         TimingData             => TmDt_WMODEA_CLKA_posedge,
         TestSignal             => WMODEA_ipd, 
         TestSignalName         => "WMODEA",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WMODEA_CLKA_posedge_posedge,
         SetupLow               => tsetup_WMODEA_CLKA_negedge_posedge,
         HoldHigh               => thold_WMODEA_CLKA_posedge_posedge,
         HoldLow                => thold_WMODEA_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     
     VitalSetupHoldCheck (
         Violation              => Tviol_DINA8_CLKA_posedge,
         TimingData             => TmDt_DINA8_CLKA_posedge,
         TestSignal             => DINA8_ipd, 
         TestSignalName         => "DINA8",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA8_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA8_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA8_CLKA_posedge_posedge,
         HoldLow                => thold_DINA8_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_DINA7_CLKA_posedge,
         TimingData             => TmDt_DINA7_CLKA_posedge,
         TestSignal             => DINA7_ipd, 
         TestSignalName         => "DINA7",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA7_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA7_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA7_CLKA_posedge_posedge,
         HoldLow                => thold_DINA7_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_DINA6_CLKA_posedge,
         TimingData             => TmDt_DINA6_CLKA_posedge,
         TestSignal             => DINA6_ipd, 
         TestSignalName         => "DINA6",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA6_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA6_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA6_CLKA_posedge_posedge,
         HoldLow                => thold_DINA6_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINA5_CLKA_posedge,
         TimingData             => TmDt_DINA5_CLKA_posedge,
         TestSignal             => DINA5_ipd, 
         TestSignalName         => "DINA5",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA5_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA5_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA5_CLKA_posedge_posedge,
         HoldLow                => thold_DINA5_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINA4_CLKA_posedge,
         TimingData             => TmDt_DINA4_CLKA_posedge,
         TestSignal             => DINA4_ipd, 
         TestSignalName         => "DINA4",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA4_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA4_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA4_CLKA_posedge_posedge,
         HoldLow                => thold_DINA4_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINA3_CLKA_posedge,
         TimingData             => TmDt_DINA3_CLKA_posedge,
         TestSignal             => DINA3_ipd, 
         TestSignalName         => "DINA3",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA3_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA3_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA3_CLKA_posedge_posedge,
         HoldLow                => thold_DINA3_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINA2_CLKA_posedge,
         TimingData             => TmDt_DINA2_CLKA_posedge,
         TestSignal             => DINA2_ipd, 
         TestSignalName         => "DINA2",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA2_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA2_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA2_CLKA_posedge_posedge,
         HoldLow                => thold_DINA2_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_DINA1_CLKA_posedge,
         TimingData             => TmDt_DINA1_CLKA_posedge,
         TestSignal             => DINA1_ipd, 
         TestSignalName         => "DINA1",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA1_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA1_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA1_CLKA_posedge_posedge,
         HoldLow                => thold_DINA1_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINA0_CLKA_posedge,
         TimingData             => TmDt_DINA0_CLKA_posedge,
         TestSignal             => DINA0_ipd, 
         TestSignalName         => "DINA0",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINA0_CLKA_posedge_posedge,
         SetupLow               => tsetup_DINA0_CLKA_negedge_posedge,
         HoldHigh               => thold_DINA0_CLKA_posedge_posedge,
         HoldLow                => thold_DINA0_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')  and
                                    (TO_X01(WENA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB8_CLKB_posedge,
         TimingData             => TmDt_DINB8_CLKB_posedge,
         TestSignal             => DINB8_ipd, 
         TestSignalName         => "DINB8",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB8_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB8_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB8_CLKB_posedge_posedge,
         HoldLow                => thold_DINB8_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB7_CLKB_posedge,
         TimingData             => TmDt_DINB7_CLKB_posedge,
         TestSignal             => DINB7_ipd, 
         TestSignalName         => "DINB7",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB7_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB7_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB7_CLKB_posedge_posedge,
         HoldLow                => thold_DINB7_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB6_CLKB_posedge,
         TimingData             => TmDt_DINB6_CLKB_posedge,
         TestSignal             => DINB6_ipd, 
         TestSignalName         => "DINB6",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB6_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB6_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB6_CLKB_posedge_posedge,
         HoldLow                => thold_DINB6_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
     
     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB5_CLKB_posedge,
         TimingData             => TmDt_DINB5_CLKB_posedge,
         TestSignal             => DINB5_ipd, 
         TestSignalName         => "DINB5",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB5_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB5_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB5_CLKB_posedge_posedge,
         HoldLow                => thold_DINB5_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB4_CLKB_posedge,
         TimingData             => TmDt_DINB4_CLKB_posedge,
         TestSignal             => DINB4_ipd, 
         TestSignalName         => "DINB4",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB4_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB4_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB4_CLKB_posedge_posedge,
         HoldLow                => thold_DINB4_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB3_CLKB_posedge,
         TimingData             => TmDt_DINB3_CLKB_posedge,
         TestSignal             => DINB3_ipd, 
         TestSignalName         => "DINB3",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB3_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB3_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB3_CLKB_posedge_posedge,
         HoldLow                => thold_DINB3_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_DINB2_CLKB_posedge,
         TimingData             => TmDt_DINB2_CLKB_posedge,
         TestSignal             => DINB2_ipd, 
         TestSignalName         => "DINB2",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB2_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB2_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB2_CLKB_posedge_posedge,
         HoldLow                => thold_DINB2_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB1_CLKB_posedge,
         TimingData             => TmDt_DINB1_CLKB_posedge,
         TestSignal             => DINB1_ipd, 
         TestSignalName         => "DINB1",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB1_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB1_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB1_CLKB_posedge_posedge,
         HoldLow                => thold_DINB1_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_DINB0_CLKB_posedge,
         TimingData             => TmDt_DINB0_CLKB_posedge,
         TestSignal             => DINB0_ipd, 
         TestSignalName         => "DINB0",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_DINB0_CLKB_posedge_posedge,
         SetupLow               => tsetup_DINB0_CLKB_negedge_posedge,
         HoldHigh               => thold_DINB0_CLKB_posedge_posedge,
         HoldLow                => thold_DINB0_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')  and
                                    (TO_X01(WENB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB11_CLKB_posedge,
         TimingData             => TmDt_ADDRB11_CLKB_posedge,
         TestSignal             => ADDRB11_ipd, 
         TestSignalName         => "ADDRB11",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB11_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB11_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB11_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB11_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB10_CLKB_posedge,
         TimingData             => TmDt_ADDRB10_CLKB_posedge,
         TestSignal             => ADDRB10_ipd, 
         TestSignalName         => "ADDRB10",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB10_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB10_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB10_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB10_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB9_CLKB_posedge,
         TimingData             => TmDt_ADDRB9_CLKB_posedge,
         TestSignal             => ADDRB9_ipd, 
         TestSignalName         => "ADDRB9",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB9_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB9_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB9_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB9_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB8_CLKB_posedge,
         TimingData             => TmDt_ADDRB8_CLKB_posedge,
         TestSignal             => ADDRB8_ipd, 
         TestSignalName         => "ADDRB8",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB8_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB8_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB8_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB8_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB7_CLKB_posedge,
         TimingData             => TmDt_ADDRB7_CLKB_posedge,
         TestSignal             => ADDRB7_ipd, 
         TestSignalName         => "ADDRB7",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB7_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB7_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB7_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB7_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB6_CLKB_posedge,
         TimingData             => TmDt_ADDRB6_CLKB_posedge,
         TestSignal             => ADDRB6_ipd, 
         TestSignalName         => "ADDRB6",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB6_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB6_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB6_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB6_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB5_CLKB_posedge,
         TimingData             => TmDt_ADDRB5_CLKB_posedge,
         TestSignal             => ADDRB5_ipd, 
         TestSignalName         => "ADDRB5",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB5_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB5_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB5_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB5_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRB4_CLKB_posedge,
         TimingData             => TmDt_ADDRB4_CLKB_posedge,
         TestSignal             => ADDRB4_ipd, 
         TestSignalName         => "ADDRB4",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB4_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB4_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB4_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB4_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRB3_CLKB_posedge,
         TimingData             => TmDt_ADDRB3_CLKB_posedge,
         TestSignal             => ADDRB3_ipd, 
         TestSignalName         => "ADDRB3",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB3_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB3_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB3_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB3_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRB2_CLKB_posedge,
         TimingData             => TmDt_ADDRB2_CLKB_posedge,
         TestSignal             => ADDRB2_ipd, 
         TestSignalName         => "ADDRB2",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB2_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB2_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB2_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB2_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB1_CLKB_posedge,
         TimingData             => TmDt_ADDRB1_CLKB_posedge,
         TestSignal             => ADDRB1_ipd, 
         TestSignalName         => "ADDRB1",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB1_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB1_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB1_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB1_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRB0_CLKB_posedge,
         TimingData             => TmDt_ADDRB0_CLKB_posedge,
         TestSignal             => ADDRB0_ipd, 
         TestSignalName         => "ADDRB0",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKB_ipd,
         RefSignalName          => "CLKB",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRB0_CLKB_posedge_posedge,
         SetupLow               => tsetup_ADDRB0_CLKB_negedge_posedge,
         HoldHigh               => thold_ADDRB0_CLKB_posedge_posedge,
         HoldLow                => thold_ADDRB0_CLKB_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA0_CLKA_posedge,
         TimingData             => TmDt_ADDRA0_CLKA_posedge,
         TestSignal             => ADDRA0_ipd, 
         TestSignalName         => "ADDRA0",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA0_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA0_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA0_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA0_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA1_CLKA_posedge,
         TimingData             => TmDt_ADDRA1_CLKA_posedge,
         TestSignal             => ADDRA1_ipd, 
         TestSignalName         => "ADDRA1",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA1_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA1_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA1_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA1_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA2_CLKA_posedge,
         TimingData             => TmDt_ADDRA2_CLKA_posedge,
         TestSignal             => ADDRA2_ipd, 
         TestSignalName         => "ADDRA2",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA2_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA2_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA2_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA2_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRA3_CLKA_posedge,
         TimingData             => TmDt_ADDRA3_CLKA_posedge,
         TestSignal             => ADDRA3_ipd, 
         TestSignalName         => "ADDRA3",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA3_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA3_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA3_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA3_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRA4_CLKA_posedge,
         TimingData             => TmDt_ADDRA4_CLKA_posedge,
         TestSignal             => ADDRA4_ipd, 
         TestSignalName         => "ADDRA4",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA4_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA4_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA4_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA4_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA5_CLKA_posedge,
         TimingData             => TmDt_ADDRA5_CLKA_posedge,
         TestSignal             => ADDRA5_ipd, 
         TestSignalName         => "ADDRA5",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA5_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA5_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA5_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA5_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA6_CLKA_posedge,
         TimingData             => TmDt_ADDRA6_CLKA_posedge,
         TestSignal             => ADDRA6_ipd, 
         TestSignalName         => "ADDRA6",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA6_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA6_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA6_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA6_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA7_CLKA_posedge,
         TimingData             => TmDt_ADDRA7_CLKA_posedge,
         TestSignal             => ADDRA7_ipd, 
         TestSignalName         => "ADDRA7",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA7_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA7_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA7_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA7_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA8_CLKA_posedge,
         TimingData             => TmDt_ADDRA8_CLKA_posedge,
         TestSignal             => ADDRA8_ipd, 
         TestSignalName         => "ADDRA8",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA8_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA8_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA8_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA8_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA9_CLKA_posedge,
         TimingData             => TmDt_ADDRA9_CLKA_posedge,
         TestSignal             => ADDRA9_ipd, 
         TestSignalName         => "ADDRA9",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA9_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA9_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA9_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA9_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck (
         Violation              => Tviol_ADDRA10_CLKA_posedge,
         TimingData             => TmDt_ADDRA10_CLKA_posedge,
         TestSignal             => ADDRA10_ipd, 
         TestSignalName         => "ADDRA10",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA10_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA10_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA10_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA10_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_ADDRA11_CLKA_posedge,
         TimingData             => TmDt_ADDRA11_CLKA_posedge,
         TestSignal             => ADDRA11_ipd, 
         TestSignalName         => "ADDRA11",
         TestDelay              => 0.0 ns,
         RefSignal              => CLKA_ipd,
         RefSignalName          => "CLKA",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_ADDRA11_CLKA_posedge_posedge,
         SetupLow               => tsetup_ADDRA11_CLKA_negedge_posedge,
         HoldHigh               => thold_ADDRA11_CLKA_posedge_posedge,
         HoldLow                => thold_ADDRA11_CLKA_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

    --  Period of CLKA
     VitalPeriodPulseCheck ( 
         Violation              => Pviol_CLKA,
         PeriodData             => PeriodData_CLKA,
         TestSignal             => CLKA_ipd, 
         TestSignalName         => "CLKA",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => tpw_CLKA_posedge,
         PulseWidthLow          => tpw_CLKA_negedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKA_ipd) = '0')),
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

    --  Period of CLKB
     VitalPeriodPulseCheck ( 
         Violation              => Pviol_CLKB,
         PeriodData             => PeriodData_CLKB,
         TestSignal             => CLKB_ipd, 
         TestSignalName         => "CLKB",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => tpw_CLKB_posedge,
         PulseWidthLow          => tpw_CLKB_negedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and
                                    (TO_X01(BLKB_ipd) = '0')),
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

    --  Period of RESET
     VitalPeriodPulseCheck ( 
         Violation              => Pviol_RESET,
         PeriodData             => PeriodData_RESET,
         TestSignal             => RESET_ipd, 
         TestSignalName         => "RESET",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => 0.0 ns,
         PulseWidthLow          => tpw_RESET_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/RAM4K9",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  end if;


  -- Calculate widthA integer value
  if ( WIDTHA1_ipd'event or WIDTHA0_ipd'event ) then
      if ((TO_X01(WIDTHA1_ipd) ='0')    and (TO_X01(WIDTHA0_ipd) ='0')) then
        widthA  := 1;
        WDA_INT := 0;
      elsif ((TO_X01(WIDTHA1_ipd) ='0') and (TO_X01(WIDTHA0_ipd) ='1')) then
        widthA  := 2;
        WDA_INT := 1;
      elsif ((TO_X01(WIDTHA1_ipd) ='1') and (TO_X01(WIDTHA0_ipd) ='0')) then
        widthA  := 4;
        WDA_INT := 2;
      elsif ((TO_X01(WIDTHA1_ipd) ='1') and (TO_X01(WIDTHA0_ipd) ='1')) then
        widthA  := 9;
        WDA_INT := 3;
      else
        widthA  := -1;
        WDA_INT := -1;
      end if;
  end if;

  -- Calculate widthB integer value
  if ( WIDTHB1_ipd'event or WIDTHB0_ipd'event ) then
      if ((TO_X01(WIDTHB1_ipd) ='0')    and (TO_X01(WIDTHB0_ipd) ='0')) then
        widthB  := 1;
        WDB_INT := 0;
      elsif ((TO_X01(WIDTHB1_ipd) ='0') and (TO_X01(WIDTHB0_ipd) ='1')) then
        widthB  := 2;
        WDB_INT := 1;
      elsif ((TO_X01(WIDTHB1_ipd) ='1') and (TO_X01(WIDTHB0_ipd) ='0')) then
        widthB  := 4;
        WDB_INT := 2;
      elsif ((TO_X01(WIDTHB1_ipd) ='1') and (TO_X01(WIDTHB0_ipd) ='1')) then
        widthB  := 9;
        WDB_INT := 3;
      else
        widthB  := -1;
        WDB_INT := -1;
      end if;
  end if;


  -----------------------------------------------------------
  --    Check if address out of range for specified width  --
  -----------------------------------------------------------
  
  if (TO_X01(RESET_ipd) = '1' and TO_X01(BLKA_delayed) = '0') then
    if (CLKA_ipd'event and TO_X01(CLKA_ipd) = '1') then

      WENA_lat := WENA_ipd;

      -- Calculate the integer address value

      ADDRA := (INT(ADDRA11_delayed)*2048) + (INT(ADDRA10_delayed)*1024) +
               (INT(ADDRA9_delayed)*512)   + (INT(ADDRA8_delayed)*256)   +
               (INT(ADDRA7_delayed)*128)   + (INT(ADDRA6_delayed)*64)    +
               (INT(ADDRA5_delayed)*32)    + (INT(ADDRA4_delayed)*16)    +
               (INT(ADDRA3_delayed)*8)     + (INT(ADDRA2_delayed)*4)     +
               (INT(ADDRA1_delayed)*2)     + (INT(ADDRA0_delayed)*1);

      if (ADDRA < 0) then
        ADDRA_VALID := 0;
      else
        ADDRA_VALID := 1;
      end if;

      if (widthA = 1 and ADDRA >= 4096) then
        ADDRA_VALID := 0;
      elsif (widthA = 2 and ADDRA >= 2048) then
        ADDRA_VALID := 0;
      elsif (widthA = 4 and ADDRA >= 1024) then
        ADDRA_VALID := 0;
      elsif (widthA = 9 and ADDRA >= 512) then
        ADDRA_VALID := 0;
      end if;

      if ( WARNING_MSGS_ON ) then
        assert (widthA /= 1 or (ADDRA < 4096 and ADDRA >= 0) )
          report "Illegal address on port A, should be between 0 & 4095."
          severity Warning;

        assert (widthA /= 2 or (ADDRA < 2048 and ADDRA >= 0) )
          report "Illegal address on port A, should be between 0 & 2047."
          severity Warning;

        assert (widthA /= 4 or (ADDRA < 1024 and ADDRA >= 0) )
          report "Illegal address on port A, should be between 0 & 1023."
          severity Warning;

        assert (widthA /= 9 or (ADDRA < 512 and ADDRA >= 0) )
          report "Illegal address on port A, should be between 0 & 511."
          severity Warning;
      end if;

    end if;
  end if;
  
  if (TO_X01(RESET_ipd) = '1' and TO_X01(BLKB_delayed) = '0') then
    if (CLKB_ipd'event and TO_X01(CLKB_ipd) = '1') then

      WENB_lat := WENB_ipd;

      -- Calculate the integer address value

      ADDRB := (INT(ADDRB11_delayed)*2048) + (INT(ADDRB10_delayed)*1024) +
               (INT(ADDRB9_delayed)*512)   + (INT(ADDRB8_delayed)*256)   +
               (INT(ADDRB7_delayed)*128)   + (INT(ADDRB6_delayed)*64)    +
               (INT(ADDRB5_delayed)*32)    + (INT(ADDRB4_delayed)*16)    +
               (INT(ADDRB3_delayed)*8)     + (INT(ADDRB2_delayed)*4)     +
               (INT(ADDRB1_delayed)*2)     + (INT(ADDRB0_delayed)*1);

      if (ADDRB < 0) then
        ADDRB_VALID := 0;
      else
        ADDRB_VALID := 1;
      end if;

      if (widthB = 1 and ADDRB >= 4096) then
        ADDRB_VALID := 0;
      elsif (widthB = 2 and ADDRB >= 2048) then
        ADDRB_VALID := 0;
      elsif (widthB = 4 and ADDRB >= 1024) then
        ADDRB_VALID := 0;
      elsif (widthB = 9 and ADDRB >= 512) then
        ADDRB_VALID := 0;
      end if;

      if ( WARNING_MSGS_ON ) then
        assert (widthB /= 1 or (ADDRB < 4096 and ADDRB >= 0) )
          report "Illegal address on port B, should be between 0 & 4095."
          severity Warning;

        assert (widthB /= 2 or (ADDRB < 2048 and ADDRB >= 0) )
          report "Illegal address on port B, should be between 0 & 2047."
          severity Warning;

        assert (widthB /= 4 or (ADDRB < 1024 and ADDRB >= 0) )
          report "Illegal address on port B, should be between 0 & 1023."
          severity Warning;

        assert (widthB /= 9 or (ADDRB < 512 and ADDRB >= 0) )
          report "Illegal address on port B, should be between 0 & 511."
          severity Warning;
      end if;

    end if;
  end if;

  -----------------------------------------------------------
  --    RESET
  -----------------------------------------------------------

  if (TO_X01(RESET_ipd) = '0') then

        case widthA is
            when 1 =>
                        DOUTA0_zd := '0';
            when 2 =>
                        DOUTA0_zd := '0';
                        DOUTA1_zd := '0';
            when 4 =>
                        DOUTA0_zd := '0';
                        DOUTA1_zd := '0';
                        DOUTA2_zd := '0';
                        DOUTA3_zd := '0';
            when 9 =>
                        DOUTA0_zd := '0';
                        DOUTA1_zd := '0';
                        DOUTA2_zd := '0';
                        DOUTA3_zd := '0';
                        DOUTA4_zd := '0';
                        DOUTA5_zd := '0';
                        DOUTA6_zd := '0';
                        DOUTA7_zd := '0';
                        DOUTA8_zd := '0';
            when others =>
                       -- if ( WARNING_MSGS_ON ) then
                       --   assert false
                       --     report "Illegal width configuration on port A."
                       --     severity Warning;
                       -- end if;
         end case;

       case widthB is
            when 1 =>
                        DOUTB0_zd := '0';
            when 2 =>
                        DOUTB0_zd  := '0';
                        DOUTB1_zd  := '0';
            when 4 =>
                        DOUTB0_zd  := '0';
                        DOUTB1_zd  := '0';
                        DOUTB2_zd  := '0';
                        DOUTB3_zd  := '0';
            when 9 =>
                        DOUTB0_zd := '0';
                        DOUTB1_zd := '0';
                        DOUTB2_zd := '0';
                        DOUTB3_zd := '0';
                        DOUTB4_zd := '0';
                        DOUTB5_zd := '0';
                        DOUTB6_zd := '0';
                        DOUTB7_zd := '0';
                        DOUTB8_zd := '0';
            when others =>
                       -- if ( WARNING_MSGS_ON ) then
                       --   assert false
                       --     report "Illegal width configuration on port B."
                       --     severity Warning;
                       -- end if;
         end case;

     if (TO_X01(PIPEA_ipd) = '1') then
       case widthA is
            when 1 =>
                        DOUTA0_stg := '0';
            when 2 =>
                        DOUTA0_stg := '0';
                        DOUTA1_stg := '0';
            when 4 =>
                        DOUTA0_stg := '0';
                        DOUTA1_stg := '0';
                        DOUTA2_stg := '0';
                        DOUTA3_stg := '0';
            when 9 =>
                        DOUTA0_stg := '0';
                        DOUTA1_stg := '0';
                        DOUTA2_stg := '0';
                        DOUTA3_stg := '0';
                        DOUTA4_stg := '0';
                        DOUTA5_stg := '0';
                        DOUTA6_stg := '0';
                        DOUTA7_stg := '0';
                        DOUTA8_stg := '0';
            when others =>
                       -- if ( WARNING_MSGS_ON ) then
                        --  assert false
                        --    report "Illegal width configuration on port A."
                        --    severity Warning;
                       -- end if;
         end case;

      end if;
   
      if (TO_X01(PIPEB_ipd) = '1') then
         case widthB is
            when 1 =>
                        DOUTB0_stg := '0';
            when 2 =>
                        DOUTB0_stg := '0';
                        DOUTB1_stg := '0';
            when 4 =>
                        DOUTB0_stg := '0';
                        DOUTB1_stg := '0';
                        DOUTB2_stg := '0';
                        DOUTB3_stg := '0';
            when 9 =>
                        DOUTB0_stg := '0';
                        DOUTB1_stg := '0';
                        DOUTB2_stg := '0';
                        DOUTB3_stg := '0';
                        DOUTB4_stg := '0';
                        DOUTB5_stg := '0';
                        DOUTB6_stg := '0';
                        DOUTB7_stg := '0';
                        DOUTB8_stg := '0';
            when others =>
                       -- if ( WARNING_MSGS_ON ) then
                        --  assert false
                        --    report "Illegal width configuration on port B."
                        --    severity Warning;
                       -- end if;
         end case;
      end if;
  end if; -- RESET

  -----------------------------------------------------------
  --    Port B Section
  -----------------------------------------------------------

  if (TO_X01(CLKB_ipd) = 'X') then
    if (TO_X01(RESET_ipd) = '1') then
      if (TO_X01(CLKB_previous) /= 'X') then
        if ( WARNING_MSGS_ON ) then
          assert false
            report "CLKB went unknown"
            severity Warning;
        end if;
      end if;
    end if;
	
	-- Falling edge on clkB
	elsif (CLKB_ipd'event and (TO_X01(CLKB_ipd) = '0') 
                        and (TO_X01(RESET_delayed) = '1')) then
    if (TO_X01(WENB_lat) = '0') and (ADDRB_VALID = 1) then -- write mode
    	
    	CLKB_wr_fe := now;
    	
  		-- Check if Write from Port A and Write from Port B are to the same address, write data is non-deterministic
			if ( (WENA_lat = '0') and same_addr(ADDRA, ADDRB, WDA_INT, WDB_INT) and
				  	                    ((CLKA_wr_fe + TC2CWWL) > CLKB_wr_fe) ) then
				assert false
				report " Port A Write and Port B Write to same address at same time. Write data conflict. Updating memory contents at conflicting address with X"
				severity warning;

				-- function call to determine conflicting write data bits based on address and width configuration
				DINB_array := drive_data_x ( ADDRA, ADDRB, WDA_INT, WDB_INT, DINB_array );
			end if;	
				-- re-assign function return value (resolved write data bits) to DINB*_delayed variables
				DINB8_delayed := DINB_array ( 8 );
				DINB7_delayed := DINB_array ( 7 );
				DINB6_delayed := DINB_array ( 6 );
				DINB5_delayed := DINB_array ( 5 );
				DINB4_delayed := DINB_array ( 4 );
				DINB3_delayed := DINB_array ( 3 );
				DINB2_delayed := DINB_array ( 2 );
				DINB1_delayed := DINB_array ( 1 );
				DINB0_delayed := DINB_array ( 0 );
				
				case (widthB) is
						when 1 =>
											 MEM_512_9 ( (ADDRB / 8), (ADDRB mod 8) ) := DINB0_delayed;
						when 2 =>
											 MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2) ) := DINB0_delayed;
											 MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2 + 1) ) := DINB1_delayed;
						when 4 =>
											 MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4) ) := DINB0_delayed;
											 MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 1) ) := DINB1_delayed;
											 MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 2) ) := DINB2_delayed;
											 MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 3) ) := DINB3_delayed;
						when 9 =>
											 MEM_512_9( (ADDRB), 0 ) := DINB0_delayed;
											 MEM_512_9( (ADDRB), 1 ) := DINB1_delayed;
											 MEM_512_9( (ADDRB), 2 ) := DINB2_delayed;
											 MEM_512_9( (ADDRB), 3 ) := DINB3_delayed;
											 MEM_512_9( (ADDRB), 4 ) := DINB4_delayed;
											 MEM_512_9( (ADDRB), 5 ) := DINB5_delayed;
											 MEM_512_9( (ADDRB), 6 ) := DINB6_delayed;
											 MEM_512_9( (ADDRB), 7 ) := DINB7_delayed;
											 MEM_512_9( (ADDRB), 8 ) := DINB8_delayed;
						when others =>
										 if ( WARNING_MSGS_ON ) then
											 assert false
												 report "Illegal width configuration on port B."
												 severity Warning;
										 end if;
				end case;
				
		end if; -- write mode
	
  elsif (CLKB_ipd'event and (TO_X01(CLKB_ipd) = '1') 
                        and (TO_X01(RESET_delayed) = '1')) then
	-- positive clk edge
    if (TO_X01(PIPEB_delayed) = '1') then -- pipelining on
      case (widthB) is
        when 1 => 
                   DOUTB0_zd   := DOUTB0_stg;
        when 2 => 
                   DOUTB0_zd   := DOUTB0_stg;
                   DOUTB1_zd   := DOUTB1_stg;
        when 4 => 
                   DOUTB0_zd   := DOUTB0_stg;
                   DOUTB1_zd   := DOUTB1_stg;
                   DOUTB2_zd   := DOUTB2_stg;
                   DOUTB3_zd   := DOUTB3_stg;
        when 9 =>  
                   DOUTB0_zd   := DOUTB0_stg;
                   DOUTB1_zd   := DOUTB1_stg;
                   DOUTB2_zd   := DOUTB2_stg;
                   DOUTB3_zd   := DOUTB3_stg;
                   DOUTB4_zd   := DOUTB4_stg;
                   DOUTB5_zd   := DOUTB5_stg;
                   DOUTB6_zd   := DOUTB6_stg;
                   DOUTB7_zd   := DOUTB7_stg;
                   DOUTB8_zd   := DOUTB8_stg;
        when others => 
                   if ( WARNING_MSGS_ON ) then
                     assert false
                       report "Illegal width configuration on port B."
                       severity Warning;
                   end if;
       end case;
    elsif (TO_X01(PIPEB_delayed) = 'X') then 
      if ( WARNING_MSGS_ON ) then
        assert false
          report "PIPEB unknown."
          severity Warning;
      end if;
      DOUTB0_zd   := 'X';
      DOUTB1_zd   := 'X';
      DOUTB2_zd   := 'X';
      DOUTB3_zd   := 'X';
      DOUTB4_zd   := 'X';
      DOUTB5_zd   := 'X';
      DOUTB6_zd   := 'X';
      DOUTB7_zd   := 'X';
      DOUTB8_zd   := 'X';
    end if; 

    if (TO_X01(BLKB_delayed) = '0') then
      if (TO_X01(WENB_delayed) ='1') and (ADDRB_VALID = 1) then -- Read mode

        CLKB_rd_re := now;

        if (TO_X01(PIPEB_delayed) = '0') then -- no pipeline
          
          -- Check if Write from Port A and Read from Port B are to the same address, read data on Port B is driven to X
          if ( (WENA_lat = '0') and same_addr(ADDRA, ADDRB, WDA_INT, WDB_INT) and
                                               ((CLKA_wr_re + TC2CWRH) > CLKB_rd_re) ) then
            assert false
            report " Port A Write and Port B Read to same address at same time. Port B read data is unpredictable, driving read data to X."
            severity warning;

            DOUTB_array := ( DOUTB8_zd & DOUTB7_zd & DOUTB6_zd & DOUTB5_zd & DOUTB4_zd &
                                           DOUTB3_zd & DOUTB2_zd & DOUTB1_zd & DOUTB0_zd );
            DOUTB_array := drive_data_x ( ADDRA, ADDRB, WDA_INT, WDB_INT, DOUTB_array );
            DOUTB8_zd := DOUTB_array ( 8 );
            DOUTB7_zd := DOUTB_array ( 7 );
            DOUTB6_zd := DOUTB_array ( 6 );
            DOUTB5_zd := DOUTB_array ( 5 );
            DOUTB4_zd := DOUTB_array ( 4 );
            DOUTB3_zd := DOUTB_array ( 3 );
            DOUTB2_zd := DOUTB_array ( 2 );
            DOUTB1_zd := DOUTB_array ( 1 );
            DOUTB0_zd := DOUTB_array ( 0 );
          else					
						case (widthB) is
	            when 1 =>
	                        DOUTB0_zd := MEM_512_9( (ADDRB / 8), (ADDRB mod 8) );
	            when 2 =>
	                        DOUTB0_zd := MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2) );
	                        DOUTB1_zd := MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2 + 1) );

	            when 4 =>
	                        DOUTB0_zd := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4) );
	                        DOUTB1_zd := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 1) );
	                        DOUTB2_zd := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 2) );
	                        DOUTB3_zd := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 3) );
	            when 9 =>
	                        DOUTB0_zd := MEM_512_9( (ADDRB), 0 );
	                        DOUTB1_zd := MEM_512_9( (ADDRB), 1 );
	                        DOUTB2_zd := MEM_512_9( (ADDRB), 2 );
	                        DOUTB3_zd := MEM_512_9( (ADDRB), 3 );
	                        DOUTB4_zd := MEM_512_9( (ADDRB), 4 );
	                        DOUTB5_zd := MEM_512_9( (ADDRB), 5 );
	                        DOUTB6_zd := MEM_512_9( (ADDRB), 6 );
	                        DOUTB7_zd := MEM_512_9( (ADDRB), 7 );
	                        DOUTB8_zd := MEM_512_9( (ADDRB), 8 );

	            when others =>
	                        if ( WARNING_MSGS_ON ) then
	                          assert false
	                            report "Illegal width configuration on port B."
	                            severity Warning;
	                        end if;
	          end case;
					end if;
        elsif (TO_X01(PIPEB_delayed) = '1') then -- pipelining on
          -- Check if Write from Port A and Read from Port B are to the same address, read data on Port B is driven to X
          if ( (WENA_lat = '0') and same_addr(ADDRA, ADDRB, WDA_INT, WDB_INT) and
                                               ((CLKA_wr_re + TC2CWRH) > CLKB_rd_re) ) then
						assert false
						report " Port A Write and Port B Read to same address at same time. Port B read data is unpredictable, driving read data to X. Updating memory contents at conflicting address with X"
						severity warning;

            DOUTB_array := ( DOUTB8_stg & DOUTB7_stg & DOUTB6_stg & DOUTB5_stg & DOUTB4_stg &
                                            DOUTB3_stg & DOUTB2_stg & DOUTB1_stg & DOUTB0_stg );
            DOUTB_array := drive_data_x ( ADDRA, ADDRB, WDA_INT, WDB_INT, DOUTB_array );
            DOUTB8_stg := DOUTB_array ( 8 );
            DOUTB7_stg := DOUTB_array ( 7 );
            DOUTB6_stg := DOUTB_array ( 6 );
            DOUTB5_stg := DOUTB_array ( 5 );
            DOUTB4_stg := DOUTB_array ( 4 );
            DOUTB3_stg := DOUTB_array ( 3 );
            DOUTB2_stg := DOUTB_array ( 2 );
            DOUTB1_stg := DOUTB_array ( 1 );
            DOUTB0_stg := DOUTB_array ( 0 );
          else
						case (widthB) is
	            when 1 =>
	                        DOUTB0_stg := MEM_512_9( (ADDRB / 8), (ADDRB mod 8) );
	            when 2 =>
	                        DOUTB0_stg := MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2) );
	                        DOUTB1_stg := MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2 + 1) );
	            when 4 =>
	                        DOUTB0_stg := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4) );
	                        DOUTB1_stg := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 1) );
	                        DOUTB2_stg := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 2) );
	                        DOUTB3_stg := MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 3) );
	            when 9 =>
	                        DOUTB0_stg := MEM_512_9( (ADDRB), 0 );
	                        DOUTB1_stg := MEM_512_9( (ADDRB), 1 );
	                        DOUTB2_stg := MEM_512_9( (ADDRB), 2 );
	                        DOUTB3_stg := MEM_512_9( (ADDRB), 3 );
	                        DOUTB4_stg := MEM_512_9( (ADDRB), 4 );
	                        DOUTB5_stg := MEM_512_9( (ADDRB), 5 );
	                        DOUTB6_stg := MEM_512_9( (ADDRB), 6 );
	                        DOUTB7_stg := MEM_512_9( (ADDRB), 7 );
	                        DOUTB8_stg := MEM_512_9( (ADDRB), 8 );

	            when others =>
	                        if ( WARNING_MSGS_ON ) then
	                          assert false
	                            report "Illegal width configuration on port B."
	                            severity Warning;
	                        end if;
	          end case;
					end if;

        else
          if ( WARNING_MSGS_ON ) then
            assert false
              report "PIPEB unknown."
              severity Warning;
          end if;
          DOUTB0_zd   := 'X';
          DOUTB1_zd   := 'X';
          DOUTB2_zd   := 'X';
          DOUTB3_zd   := 'X';
          DOUTB4_zd   := 'X';
          DOUTB5_zd   := 'X';
          DOUTB6_zd   := 'X';
          DOUTB7_zd   := 'X';
          DOUTB8_zd   := 'X';
        end if;
      elsif (TO_X01(WENB_delayed) = '0') and (ADDRB_VALID = 1) then -- Write mode

        CLKB_wr_re := now;
				DINB_array := ( DINB8_delayed & DINB7_delayed & DINB6_delayed & DINB5_delayed & DINB4_delayed &
                                            DINB3_delayed & DINB2_delayed & DINB1_delayed & DINB0_delayed );

				-- if no conflicting writes, assign write data to bypass variables, DINA*_bypass for driving onto RD if MODE=1
				DINB8_bypass := DINB8_delayed;
				DINB7_bypass := DINB7_delayed;
				DINB6_bypass := DINB6_delayed;
				DINB5_bypass := DINB5_delayed;
				DINB4_bypass := DINB4_delayed;
				DINB3_bypass := DINB3_delayed;
				DINB2_bypass := DINB2_delayed;
				DINB1_bypass := DINB1_delayed;
				DINB0_bypass := DINB0_delayed;

        -- Check if Read from Port A and Write from Port B are to the same address, write data is non-deterministic
        if ( (WENA_lat = '1') and same_addr(ADDRA, ADDRB, WDA_INT, WDB_INT) and
                                             ((CLKA_rd_re + TC2CRWH) > CLKB_wr_re) ) then
            assert false
            report " Port A Read and Port B Write to same address at same time. Port A read data is unpredictable, driving read data to X."
            severity warning;

            if (TO_X01(PIPEA_delayed) = '1') then -- pipelining on
              DOUTA_array := ( DOUTA8_stg & DOUTA7_stg & DOUTA6_stg & DOUTA5_stg & DOUTA4_stg &
                                             DOUTA3_stg & DOUTA2_stg & DOUTA1_stg & DOUTA0_stg );
              DOUTA_array := drive_data_x ( ADDRB, ADDRA, WDB_INT, WDA_INT, DOUTA_array );
              DOUTA8_stg := DOUTA_array ( 8 );
              DOUTA7_stg := DOUTA_array ( 7 );
              DOUTA6_stg := DOUTA_array ( 6 );
              DOUTA5_stg := DOUTA_array ( 5 );
              DOUTA4_stg := DOUTA_array ( 4 );
              DOUTA3_stg := DOUTA_array ( 3 );
              DOUTA2_stg := DOUTA_array ( 2 );
              DOUTA1_stg := DOUTA_array ( 1 );
              DOUTA0_stg := DOUTA_array ( 0 );
            elsif (TO_X01(PIPEA_delayed) = '0') then -- pipelining off
              DOUTA_array := ( DOUTA8_zd & DOUTA7_zd & DOUTA6_zd & DOUTA5_zd & DOUTA4_zd &
                                             DOUTA3_zd & DOUTA2_zd & DOUTA1_zd & DOUTA0_zd );
              DOUTA_array := drive_data_x ( ADDRB, ADDRA, WDB_INT, WDA_INT, DOUTA_array );
              DOUTA8_zd := DOUTA_array ( 8 );
              DOUTA7_zd := DOUTA_array ( 7 );
              DOUTA6_zd := DOUTA_array ( 6 );
              DOUTA5_zd := DOUTA_array ( 5 );
              DOUTA4_zd := DOUTA_array ( 4 );
              DOUTA3_zd := DOUTA_array ( 3 );
              DOUTA2_zd := DOUTA_array ( 2 );
              DOUTA1_zd := DOUTA_array ( 1 );
              DOUTA0_zd := DOUTA_array ( 0 );
            end if;
				end if;

        case (widthB) is
            when 1 =>
                       MEM_512_9 ( (ADDRB / 8), (ADDRB mod 8) ) := DINB0_delayed;

                       if (TO_X01(WMODEB_ipd) = '1') then
                         if (TO_X01(PIPEB_ipd) = '0') then
                           DOUTB0_zd := DINB0_bypass;
                         elsif (TO_X01(PIPEB_ipd) = '1') then
                           DOUTB0_stg := DINB0_bypass;
                         end if;
                       end if;
            when 2 =>
                       MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2) ) := DINB0_delayed;
                       MEM_512_9( (ADDRB / 4), ((ADDRB mod 4) * 2 + 1) ) := DINB1_delayed;

                       if (TO_X01(WMODEB_ipd) = '1') then
                         if (TO_X01(PIPEB_ipd) = '0') then
                           DOUTB0_zd := DINB0_bypass;
                           DOUTB1_zd := DINB1_bypass;
                         elsif (TO_X01(PIPEB_ipd) = '1') then
                           DOUTB0_stg := DINB0_bypass;
                           DOUTB1_stg := DINB1_bypass;
                         end if;
                       end if;

            when 4 =>
                       MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4) ) := DINB0_delayed;
                       MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 1) ) := DINB1_delayed;
                       MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 2) ) := DINB2_delayed;
                       MEM_512_9( (ADDRB / 2), ((ADDRB mod 2) * 4 + 3) ) := DINB3_delayed;

                       if (TO_X01(WMODEB_ipd) = '1') then
                         if (TO_X01(PIPEB_ipd) = '0') then
                           DOUTB0_zd := DINB0_bypass;
                           DOUTB1_zd := DINB1_bypass;
                           DOUTB2_zd := DINB2_bypass;
                           DOUTB3_zd := DINB3_bypass;
                         elsif (TO_X01(PIPEB_ipd) = '1') then
                           DOUTB0_stg := DINB0_bypass;
                           DOUTB1_stg := DINB1_bypass;
                           DOUTB2_stg := DINB2_bypass;
                           DOUTB3_stg := DINB3_bypass;
                         end if;
                       end if;
            when 9 =>
                       MEM_512_9( (ADDRB), 0 ) := DINB0_delayed;
                       MEM_512_9( (ADDRB), 1 ) := DINB1_delayed;
                       MEM_512_9( (ADDRB), 2 ) := DINB2_delayed;
                       MEM_512_9( (ADDRB), 3 ) := DINB3_delayed;
                       MEM_512_9( (ADDRB), 4 ) := DINB4_delayed;
                       MEM_512_9( (ADDRB), 5 ) := DINB5_delayed;
                       MEM_512_9( (ADDRB), 6 ) := DINB6_delayed;
                       MEM_512_9( (ADDRB), 7 ) := DINB7_delayed;
                       MEM_512_9( (ADDRB), 8 ) := DINB8_delayed;
 
                       if (TO_X01(WMODEB_ipd) = '1') then
                         if (TO_X01(PIPEB_ipd) = '0') then
                           DOUTB0_zd := DINB0_bypass;
                           DOUTB1_zd := DINB1_bypass;
                           DOUTB2_zd := DINB2_bypass;
                           DOUTB3_zd := DINB3_bypass;
                           DOUTB4_zd := DINB4_bypass;
                           DOUTB5_zd := DINB5_bypass;
                           DOUTB6_zd := DINB6_bypass;
                           DOUTB7_zd := DINB7_bypass;
                           DOUTB8_zd := DINB8_bypass;
                         elsif (TO_X01(PIPEB_ipd) = '1') then
                           DOUTB0_stg := DINB0_bypass;
                           DOUTB1_stg := DINB1_bypass;
                           DOUTB2_stg := DINB2_bypass;
                           DOUTB3_stg := DINB3_bypass;
                           DOUTB4_stg := DINB4_bypass;
                           DOUTB5_stg := DINB5_bypass;
                           DOUTB6_stg := DINB6_bypass;
                           DOUTB7_stg := DINB7_bypass;
                           DOUTB8_stg := DINB8_bypass;
                         end if;
                       end if;
            when others =>
                       if ( WARNING_MSGS_ON ) then
                         assert false
                           report "Illegal width configuration on port B."
                           severity Warning;
                       end if;
        end case;
      elsif (TO_X01(WENB_delayed) ='1') and (ADDRB_VALID = 0) then -- illegal read address, no read
          if ( WARNING_MSGS_ON ) then
            assert false
              report "Illegal Read Address on port B, Read Not Initiated."
              severity Warning;
          end if;
      elsif (TO_X01(WENB_delayed) ='0') and (ADDRB_VALID = 0) then -- illegal write address, no write
          if ( WARNING_MSGS_ON ) then
            assert false
              report "Illegal Write Address on port B, Write Not Initiated."
              severity Warning;
          end if;
      else
        if ( WARNING_MSGS_ON ) then
          assert false
            report "WENB unknown."
            severity Warning;
        end if;
      end if;
    elsif (TO_X01(BLKB_delayed) /= '1') then
      if ( WARNING_MSGS_ON ) then
        assert false
          report "BLKB unknown."
          severity Warning;
      end if;
    end if;
  end if;

  -----------------------------------------------------------
  --    Port A Section
  -----------------------------------------------------------

  if (TO_X01(CLKA_ipd) = 'X') then
    if (TO_X01(RESET_ipd) = '1') then
      if (TO_X01(CLKA_previous) /= 'X') then
        if ( WARNING_MSGS_ON ) then
          assert false
            report "CLKA went unknown"
            severity Warning;
        end if;
      end if;
    end if;
	
		-- Falling edge on clkA  
		elsif (CLKA_ipd'event and (TO_X01(CLKA_ipd) = '0')
													and (TO_X01(RESET_delayed) = '1')) then  
			if (TO_X01(WENA_lat) = '0') and (ADDRA_VALID = 1) then -- write mode
				CLKA_wr_fe := now;  
				-- Check if Write from Port A and Write from Port B are to the same address, write data is non-deterministic
				if ( (WENB_lat = '0') and same_addr(ADDRA, ADDRB, WDA_INT, WDB_INT) and
											((CLKB_wr_fe + TC2CWWL) > CLKA_wr_fe) ) then
					assert false
					report " Port A Write and Port B Write to same address at same time. Write data conflict. Updating memory contents at conflicting address with X"
					severity warning;

					-- function call to determine conflicting write data bits based on address and width configuration
					DINA_array := drive_data_x ( ADDRB, ADDRA, WDB_INT, WDA_INT, DINA_array );
				end if;		
					-- re-assign function return value (resolved write data bits) to DINA*_delayed variables
					DINA8_delayed := DINA_array ( 8 );
					DINA7_delayed := DINA_array ( 7 );
					DINA6_delayed := DINA_array ( 6 );
					DINA5_delayed := DINA_array ( 5 );
					DINA4_delayed := DINA_array ( 4 );
					DINA3_delayed := DINA_array ( 3 );
					DINA2_delayed := DINA_array ( 2 );
					DINA1_delayed := DINA_array ( 1 );
					DINA0_delayed := DINA_array ( 0 );
					
					
					case (widthA) is
							when 1 =>
												 MEM_512_9 ( (ADDRA / 8), (ADDRA mod 8) ) := DINA0_delayed; 
							when 2 =>
												 MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2) ) := DINA0_delayed;
												 MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2 + 1) ) := DINA1_delayed;
							when 4 =>
												 MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4) ) := DINA0_delayed;
												 MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 1) ) := DINA1_delayed;
												 MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 2) ) := DINA2_delayed;
												 MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 3) ) := DINA3_delayed;
							when 9 =>
												 MEM_512_9( (ADDRA), 0 ) := DINA0_delayed;
												 MEM_512_9( (ADDRA), 1 ) := DINA1_delayed;
												 MEM_512_9( (ADDRA), 2 ) := DINA2_delayed;
												 MEM_512_9( (ADDRA), 3 ) := DINA3_delayed;
												 MEM_512_9( (ADDRA), 4 ) := DINA4_delayed;
												 MEM_512_9( (ADDRA), 5 ) := DINA5_delayed;
												 MEM_512_9( (ADDRA), 6 ) := DINA6_delayed;
												 MEM_512_9( (ADDRA), 7 ) := DINA7_delayed;
												 MEM_512_9( (ADDRA), 8 ) := DINA8_delayed;
							when others =>
												 if ( WARNING_MSGS_ON ) then
													 assert false
														 report "Illegal width configuration on port A."
														 severity Warning;
												 end if;
					end case;
			
					
				
			end if; -- write mode
			
			
			
			
			
	
  elsif (CLKA_ipd'event and (TO_X01(CLKA_ipd) = '1')
                        and (TO_X01(RESET_delayed) = '1')) then
		-- positive clk edge
        if (TO_X01(PIPEA_delayed) = '1') then -- pipelining on
          case (widthA) is
            when 1 => 
                        DOUTA0_zd   := DOUTA0_stg;
            when 2 => 
                        DOUTA0_zd   := DOUTA0_stg;
                        DOUTA1_zd   := DOUTA1_stg;
            when 4 => 
                        DOUTA0_zd   := DOUTA0_stg;
                        DOUTA1_zd   := DOUTA1_stg;
                        DOUTA2_zd   := DOUTA2_stg;
                        DOUTA3_zd   := DOUTA3_stg;
            when 9 =>  
                        DOUTA0_zd   := DOUTA0_stg;
                        DOUTA1_zd   := DOUTA1_stg;
                        DOUTA2_zd   := DOUTA2_stg;
                        DOUTA3_zd   := DOUTA3_stg;
                        DOUTA4_zd   := DOUTA4_stg;
                        DOUTA5_zd   := DOUTA5_stg;
                        DOUTA6_zd   := DOUTA6_stg;
                        DOUTA7_zd   := DOUTA7_stg;
                        DOUTA8_zd   := DOUTA8_stg;
            when others => 
                        if ( WARNING_MSGS_ON ) then
                          assert false
                            report "Illegal width configuration on port A."
                            severity Warning;
                        end if;
          end case;
        elsif (TO_X01(PIPEA_delayed) = 'X') then
          if ( WARNING_MSGS_ON ) then
            assert false
              report "PIPEA unknown."
              severity Warning;
          end if;
          DOUTA0_zd   := 'X';
          DOUTA1_zd   := 'X';
          DOUTA2_zd   := 'X';
          DOUTA3_zd   := 'X';
          DOUTA4_zd   := 'X';
          DOUTA5_zd   := 'X';
          DOUTA6_zd   := 'X';
          DOUTA7_zd   := 'X';
          DOUTA8_zd   := 'X';
        end if; 

    if (TO_X01(BLKA_delayed) = '0') then
      if (TO_X01(WENA_delayed) = '1') and (ADDRA_VALID = 1) then -- Read mode

        CLKA_rd_re := now;

        if (TO_X01(PIPEA_delayed) = '0') then -- no pipeline
          -- Check if Write from Port B and Read from Port A are to the same address, read data on Port A is driven to X
          if ( (WENB_lat = '0') and same_addr(ADDRB, ADDRA, WDB_INT, WDA_INT) and
                                               ((CLKB_wr_re + TC2CWRH) > CLKA_rd_re) ) then
						assert false
						report " Port B Write and Port A Read to same address at same time. Port A read data is unpredictable, driving read data to X."
						severity warning;

            DOUTA_array := ( DOUTA8_zd & DOUTA7_zd & DOUTA6_zd & DOUTA5_zd & DOUTA4_zd &
                                           DOUTA3_zd & DOUTA2_zd & DOUTA1_zd & DOUTA0_zd );
            DOUTA_array := drive_data_x ( ADDRB, ADDRA, WDB_INT, WDA_INT, DOUTA_array );
            DOUTA8_zd := DOUTA_array ( 8 );
            DOUTA7_zd := DOUTA_array ( 7 );
            DOUTA6_zd := DOUTA_array ( 6 );
            DOUTA5_zd := DOUTA_array ( 5 );
            DOUTA4_zd := DOUTA_array ( 4 );
            DOUTA3_zd := DOUTA_array ( 3 );
            DOUTA2_zd := DOUTA_array ( 2 );
            DOUTA1_zd := DOUTA_array ( 1 );
            DOUTA0_zd := DOUTA_array ( 0 );
          else
						case widthA is
	            when 1 => 
	                        DOUTA0_zd := MEM_512_9( (ADDRA / 8), (ADDRA mod 8) );
	            when 2 => 
	                        DOUTA0_zd := MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2) );
	                        DOUTA1_zd := MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2 + 1) );
	            when 4 => 
	                        DOUTA0_zd := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4) );
	                        DOUTA1_zd := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 1) );
	                        DOUTA2_zd := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 2) );
	                        DOUTA3_zd := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 3) );
	            when 9 =>  
	                        DOUTA0_zd := MEM_512_9( (ADDRA), 0 );
	                        DOUTA1_zd := MEM_512_9( (ADDRA), 1 );
	                        DOUTA2_zd := MEM_512_9( (ADDRA), 2 );
	                        DOUTA3_zd := MEM_512_9( (ADDRA), 3 );
	                        DOUTA4_zd := MEM_512_9( (ADDRA), 4 );
	                        DOUTA5_zd := MEM_512_9( (ADDRA), 5 );
	                        DOUTA6_zd := MEM_512_9( (ADDRA), 6 );
	                        DOUTA7_zd := MEM_512_9( (ADDRA), 7 );
	                        DOUTA8_zd := MEM_512_9( (ADDRA), 8 );
	            when others =>
	                        if ( WARNING_MSGS_ON ) then
	                          assert false
	                            report "Illegal width configuration on port A."
	                            severity Warning;
	                        end if;
	          end case;  
					end if;

          

        elsif (TO_X01(PIPEA_delayed) = '1') then -- pipelining on
          -- Check if Write from Port B and Read from Port A are to the same address, read data on Port A is driven to X
          if ( (WENB_lat = '0') and same_addr(ADDRB, ADDRA, WDB_INT, WDA_INT) and
                                               ((CLKB_wr_re + TC2CWRH) > CLKA_rd_re) ) then
						assert false
						report " Port B Write and Port A Read to same address at same time. Port A read data is unpredictable, driving read data to X."
						severity warning;

            DOUTA_array := ( DOUTA8_stg & DOUTA7_stg & DOUTA6_stg & DOUTA5_stg & DOUTA4_stg &
                                            DOUTA3_stg & DOUTA2_stg & DOUTA1_stg & DOUTA0_stg );
            DOUTA_array := drive_data_x ( ADDRB, ADDRA, WDB_INT, WDA_INT, DOUTA_array );
            DOUTA8_stg := DOUTA_array ( 8 );
            DOUTA7_stg := DOUTA_array ( 7 );
            DOUTA6_stg := DOUTA_array ( 6 );
            DOUTA5_stg := DOUTA_array ( 5 );
            DOUTA4_stg := DOUTA_array ( 4 );
            DOUTA3_stg := DOUTA_array ( 3 );
            DOUTA2_stg := DOUTA_array ( 2 );
            DOUTA1_stg := DOUTA_array ( 1 );
            DOUTA0_stg := DOUTA_array ( 0 );
						
          else
						case (widthA) is
	            when 1 => 
	                        DOUTA0_stg := MEM_512_9( (ADDRA / 8), (ADDRA mod 8) );
	            when 2 => 
	                        DOUTA0_stg := MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2) );
	                        DOUTA1_stg := MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2 + 1) );
	            when 4 => 
	                        DOUTA0_stg := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4) );
	                        DOUTA1_stg := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 1) );
	                        DOUTA2_stg := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 2) );
	                        DOUTA3_stg := MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 3) );
	            when 9 => 
	                        DOUTA0_stg := MEM_512_9( (ADDRA), 0 );
	                        DOUTA1_stg := MEM_512_9( (ADDRA), 1 );
	                        DOUTA2_stg := MEM_512_9( (ADDRA), 2 );
	                        DOUTA3_stg := MEM_512_9( (ADDRA), 3 );
	                        DOUTA4_stg := MEM_512_9( (ADDRA), 4 );
	                        DOUTA5_stg := MEM_512_9( (ADDRA), 5 );
	                        DOUTA6_stg := MEM_512_9( (ADDRA), 6 );
	                        DOUTA7_stg := MEM_512_9( (ADDRA), 7 );
	                        DOUTA8_stg := MEM_512_9( (ADDRA), 8 );
	            when others => 
	                        if ( WARNING_MSGS_ON ) then
	                          assert false
	                            report "Illegal width configuration on port A."
	                            severity Warning;
	                        end if;
	          end case;
					end if;

        else 
          if ( WARNING_MSGS_ON ) then
            assert false
              report "PIPEA unknown."
              severity Warning;
          end if;
          DOUTA0_zd   := 'X';
          DOUTA1_zd   := 'X';
          DOUTA2_zd   := 'X';
          DOUTA3_zd   := 'X';
          DOUTA4_zd   := 'X';
          DOUTA5_zd   := 'X';
          DOUTA6_zd   := 'X';
          DOUTA7_zd   := 'X';
          DOUTA8_zd   := 'X';
        end if; 

      elsif (TO_X01(WENA_delayed) = '0') and (ADDRA_VALID = 1) then -- Write mode

        CLKA_wr_re := now;
				DINA_array := ( DINA8_delayed & DINA7_delayed & DINA6_delayed & DINA5_delayed & DINA4_delayed &
                                            DINA3_delayed & DINA2_delayed & DINA1_delayed & DINA0_delayed );

        -- if no conflicting writes, assign write data to bypass variables, DINA*_bypass for driving onto RD if MODE=1
				DINA8_bypass := DINA8_delayed;
				DINA7_bypass := DINA7_delayed; 
				DINA6_bypass := DINA6_delayed; 
				DINA5_bypass := DINA5_delayed;
				DINA4_bypass := DINA4_delayed;
				DINA3_bypass := DINA3_delayed;
				DINA2_bypass := DINA2_delayed;
				DINA1_bypass := DINA1_delayed;
				DINA0_bypass := DINA0_delayed;

        -- Check if Read from Port B and Write from Port A are to the same address, write data is non-deterministic
        if ( (WENB_lat = '1') and same_addr( ADDRB,  ADDRA, WDB_INT, WDA_INT) and
                                             ((CLKB_rd_re + TC2CRWH) > CLKA_wr_re) ) then
            assert false
              report " Port B Read and Port A Write to same address at same time. Port B read data is unpredictable, driving read data to X."
              severity warning;

            if (TO_X01(PIPEB_ipd) = '1') then -- pipelining on
              DOUTB_array := ( DOUTB8_stg & DOUTB7_stg & DOUTB6_stg & DOUTB5_stg & DOUTB4_stg &
                                           DOUTB3_stg & DOUTB2_stg & DOUTB1_stg & DOUTB0_stg );
              DOUTB_array := drive_data_x ( ADDRA, ADDRB, WDA_INT, WDB_INT, DOUTB_array );
              DOUTB8_stg := DOUTB_array ( 8 );
              DOUTB7_stg := DOUTB_array ( 7 );
              DOUTB6_stg := DOUTB_array ( 6 );
              DOUTB5_stg := DOUTB_array ( 5 );
              DOUTB4_stg := DOUTB_array ( 4 );
              DOUTB3_stg := DOUTB_array ( 3 );
              DOUTB2_stg := DOUTB_array ( 2 );
              DOUTB1_stg := DOUTB_array ( 1 );
              DOUTB0_stg := DOUTB_array ( 0 );
            elsif (TO_X01(PIPEB_ipd) = '0') then -- pipelining off
              DOUTB_array := ( DOUTB8_zd & DOUTB7_zd & DOUTB6_zd & DOUTB5_zd & DOUTB4_zd &
                                             DOUTB3_zd & DOUTB2_zd & DOUTB1_zd & DOUTB0_zd );
              DOUTB_array := drive_data_x ( ADDRA, ADDRB, WDA_INT, WDB_INT, DOUTB_array );
              DOUTB8_zd := DOUTB_array ( 8 );
              DOUTB7_zd := DOUTB_array ( 7 );
              DOUTB6_zd := DOUTB_array ( 6 );
              DOUTB5_zd := DOUTB_array ( 5 );
              DOUTB4_zd := DOUTB_array ( 4 );
              DOUTB3_zd := DOUTB_array ( 3 );
              DOUTB2_zd := DOUTB_array ( 2 );
              DOUTB1_zd := DOUTB_array ( 1 );
              DOUTB0_zd := DOUTB_array ( 0 );
            end if;
				end if;

        case (widthA) is
            when 1 =>
                       MEM_512_9 ( (ADDRA / 8), (ADDRA mod 8) ) := DINA0_delayed; 

                       if (TO_X01(WMODEA_ipd) = '1') then 
                         if (TO_X01(PIPEA_ipd) = '0') then 
                           DOUTA0_zd := DINA0_bypass;
                         elsif (TO_X01(PIPEA_ipd) = '1') then 
                           DOUTA0_stg := DINA0_bypass;
                         end if;
                       end if;
            when 2 =>
                       MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2) ) := DINA0_delayed;
                       MEM_512_9( (ADDRA / 4), ((ADDRA mod 4) * 2 + 1) ) := DINA1_delayed;
 
                       if (TO_X01(WMODEA_ipd) = '1') then 
                         if (TO_X01(PIPEA_ipd) = '0') then 
                           DOUTA0_zd := DINA0_bypass;
                           DOUTA1_zd := DINA1_bypass;
                         elsif (TO_X01(PIPEA_ipd) = '1') then 
                           DOUTA0_stg := DINA0_bypass;
                           DOUTA1_stg := DINA1_bypass;
                         end if;
                       end if;
            when 4 =>
                       MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4) ) := DINA0_delayed;
                       MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 1) ) := DINA1_delayed;
                       MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 2) ) := DINA2_delayed;
                       MEM_512_9( (ADDRA / 2), ((ADDRA mod 2) * 4 + 3) ) := DINA3_delayed;

                       if (TO_X01(WMODEA_ipd) = '1') then 
                         if (TO_X01(PIPEA_ipd) = '0') then 
                           DOUTA0_zd := DINA0_bypass;
                           DOUTA1_zd := DINA1_bypass;
                           DOUTA2_zd := DINA2_bypass;
                           DOUTA3_zd := DINA3_bypass;
                         elsif (TO_X01(PIPEA_ipd) = '1') then 
                           DOUTA0_stg := DINA0_bypass;
                           DOUTA1_stg := DINA1_bypass;
                           DOUTA2_stg := DINA2_bypass;
                           DOUTA3_stg := DINA3_bypass;
                         end if;
                       end if;
            when 9 =>
                       MEM_512_9( (ADDRA), 0 ) := DINA0_delayed;
                       MEM_512_9( (ADDRA), 1 ) := DINA1_delayed;
                       MEM_512_9( (ADDRA), 2 ) := DINA2_delayed;
                       MEM_512_9( (ADDRA), 3 ) := DINA3_delayed;
                       MEM_512_9( (ADDRA), 4 ) := DINA4_delayed;
                       MEM_512_9( (ADDRA), 5 ) := DINA5_delayed;
                       MEM_512_9( (ADDRA), 6 ) := DINA6_delayed;
                       MEM_512_9( (ADDRA), 7 ) := DINA7_delayed;
                       MEM_512_9( (ADDRA), 8 ) := DINA8_delayed;
                       
                       if (TO_X01(WMODEA_ipd) = '1') then 
                         if (TO_X01(PIPEA_ipd) = '0') then 
                           DOUTA0_zd := DINA0_bypass;
                           DOUTA1_zd := DINA1_bypass;
                           DOUTA2_zd := DINA2_bypass;
                           DOUTA3_zd := DINA3_bypass;
                           DOUTA4_zd := DINA4_bypass;
                           DOUTA5_zd := DINA5_bypass;
                           DOUTA6_zd := DINA6_bypass;
                           DOUTA7_zd := DINA7_bypass;
                           DOUTA8_zd := DINA8_bypass;
                         elsif(TO_X01(PIPEA_ipd) = '1') then 
                           DOUTA0_stg := DINA0_bypass;
                           DOUTA1_stg := DINA1_bypass;
                           DOUTA2_stg := DINA2_bypass;
                           DOUTA3_stg := DINA3_bypass;
                           DOUTA4_stg := DINA4_bypass;
                           DOUTA5_stg := DINA5_bypass;
                           DOUTA6_stg := DINA6_bypass;
                           DOUTA7_stg := DINA7_bypass;
                           DOUTA8_stg := DINA8_bypass;
                         end if;
                       end if;
            when others =>
                       if ( WARNING_MSGS_ON ) then
                         assert false
                           report "Illegal width configuration on port A."
                           severity Warning;
                       end if;
        end case;
      elsif (TO_X01(WENA_delayed) ='1') and (ADDRA_VALID = 0) then -- illegal read address, no read
          if ( WARNING_MSGS_ON ) then
            assert false
              report "Illegal Read Address on port A, Read Not Initiated."
              severity Warning;
          end if;
      elsif (TO_X01(WENA_delayed) ='0') and (ADDRA_VALID = 0) then -- illegal write address, no write
          if ( WARNING_MSGS_ON ) then
            assert false
              report "Illegal Write Address on port A, Write Not Initiated."
              severity Warning;
          end if;
      else
        if ( WARNING_MSGS_ON ) then
          assert false
            report "WENA unknown."
            severity Warning;
        end if;
      end if; 
    elsif (TO_X01(BLKA_delayed) /= '1') then
      if ( WARNING_MSGS_ON ) then
        assert false
          report "BLKA unknown."
          severity Warning;
      end if;
    end if; 
  end if;

  -----------------------------------------------------------
  --    Delayed Signals Section
  -----------------------------------------------------------

  if (CLKA'event) then
    CLKA_previous := CLKA_ipd;
  end if;

  if (CLKB'event) then
    CLKB_previous := CLKB_ipd;
  end if;
   
  WENA_delayed      := WENA_ipd;
  WENB_delayed      := WENB_ipd;
  PIPEA_delayed     := PIPEA_ipd;
  PIPEB_delayed     := PIPEB_ipd;
  RESET_delayed     := RESET_ipd;

  ADDRA11_delayed   := ADDRA11_ipd;
  ADDRA10_delayed   := ADDRA10_ipd;
  ADDRA9_delayed    := ADDRA9_ipd;
  ADDRA8_delayed    := ADDRA8_ipd;
  ADDRA7_delayed    := ADDRA7_ipd;
  ADDRA6_delayed    := ADDRA6_ipd;
  ADDRA5_delayed    := ADDRA5_ipd;
  ADDRA4_delayed    := ADDRA4_ipd;
  ADDRA3_delayed    := ADDRA3_ipd;
  ADDRA2_delayed    := ADDRA2_ipd;
  ADDRA1_delayed    := ADDRA1_ipd;
  ADDRA0_delayed    := ADDRA0_ipd;

  ADDRB11_delayed   := ADDRB11_ipd;
  ADDRB10_delayed   := ADDRB10_ipd;
  ADDRB9_delayed    := ADDRB9_ipd;
  ADDRB8_delayed    := ADDRB8_ipd;
  ADDRB7_delayed    := ADDRB7_ipd;
  ADDRB6_delayed    := ADDRB6_ipd;
  ADDRB5_delayed    := ADDRB5_ipd;
  ADDRB4_delayed    := ADDRB4_ipd;
  ADDRB3_delayed    := ADDRB3_ipd;
  ADDRB2_delayed    := ADDRB2_ipd;
  ADDRB1_delayed    := ADDRB1_ipd;
  ADDRB0_delayed    := ADDRB0_ipd;

  DINA8_delayed     := DINA8_ipd;
  DINA7_delayed     := DINA7_ipd;
  DINA6_delayed     := DINA6_ipd;
  DINA5_delayed     := DINA5_ipd;
  DINA4_delayed     := DINA4_ipd;
  DINA3_delayed     := DINA3_ipd;
  DINA2_delayed     := DINA2_ipd;
  DINA1_delayed     := DINA1_ipd;
  DINA0_delayed     := DINA0_ipd;

  DINB8_delayed     := DINB8_ipd;
  DINB7_delayed     := DINB7_ipd;
  DINB6_delayed     := DINB6_ipd;
  DINB5_delayed     := DINB5_ipd;
  DINB4_delayed     := DINB4_ipd;
  DINB3_delayed     := DINB3_ipd;
  DINB2_delayed     := DINB2_ipd;
  DINB1_delayed     := DINB1_ipd;
  DINB0_delayed     := DINB0_ipd;

  BLKA_delayed      := BLKA_ipd;
  BLKB_delayed      := BLKB_ipd;


  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

  VitalPathDelay01Z (
        OutSignal     => DOUTA0,
        GlitchData    => DOUTA0_GlitchData,
        OutSignalName => "DOUTA0",
        OutTemp       => DOUTA0_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA0), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA0), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTA1,
        GlitchData    => DOUTA1_GlitchData,
        OutSignalName => "DOUTA1",
        OutTemp       => DOUTA1_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA1), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA1), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


     
  VitalPathDelay01Z (
        OutSignal     => DOUTA2,
        GlitchData    => DOUTA2_GlitchData,
        OutSignalName => "DOUTA2",
        OutTemp       => DOUTA2_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA2), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA2), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTA3,
        GlitchData    => DOUTA3_GlitchData,
        OutSignalName => "DOUTA3",
        OutTemp       => DOUTA3_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA3), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA3), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

     
  VitalPathDelay01Z (
        OutSignal     => DOUTA4,
        GlitchData    => DOUTA4_GlitchData,
        OutSignalName => "DOUTA4",
        OutTemp       => DOUTA4_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA4), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA4), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTA5,
        GlitchData    => DOUTA5_GlitchData,
        OutSignalName => "DOUTA5",
        OutTemp       => DOUTA5_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA5), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA5), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


  VitalPathDelay01Z (
        OutSignal     => DOUTA6,
        GlitchData    => DOUTA6_GlitchData,
        OutSignalName => "DOUTA6",
        OutTemp       => DOUTA6_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA6), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA6), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

     
  VitalPathDelay01Z (
        OutSignal     => DOUTA7,
        GlitchData    => DOUTA7_GlitchData,
        OutSignalName => "DOUTA7",
        OutTemp       => DOUTA7_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA7), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA7), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTA8,
        GlitchData    => DOUTA8_GlitchData,
        OutSignalName => "DOUTA8",
        OutTemp       => DOUTA8_zd,
        Paths         => (0 => (CLKA_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKA_DOUTA8), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTA8), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


  VitalPathDelay01Z (
        OutSignal     => DOUTB0,
        GlitchData    => DOUTB0_GlitchData,
        OutSignalName => "DOUTB0",
        OutTemp       => DOUTB0_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB0), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB0), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


  VitalPathDelay01Z (
        OutSignal     => DOUTB1,
        GlitchData    => DOUTB1_GlitchData,
        OutSignalName => "DOUTB1",
        OutTemp       => DOUTB1_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB1), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB1), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTB2,
        GlitchData    => DOUTB2_GlitchData,
        OutSignalName => "DOUTB2",
        OutTemp       => DOUTB2_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB2), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB2), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTB3,
        GlitchData    => DOUTB3_GlitchData,
        OutSignalName => "DOUTB3",
        OutTemp       => DOUTB3_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB3), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB3), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


  VitalPathDelay01Z (
        OutSignal     => DOUTB4,
        GlitchData    => DOUTB4_GlitchData,
        OutSignalName => "DOUTB4",
        OutTemp       => DOUTB4_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB4), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB4), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTB5,
        GlitchData    => DOUTB5_GlitchData,
        OutSignalName => "DOUTB5",
        OutTemp       => DOUTB5_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB5), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB5), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


  VitalPathDelay01Z (
        OutSignal     => DOUTB6,
        GlitchData    => DOUTB6_GlitchData,
        OutSignalName => "DOUTB6",
        OutTemp       => DOUTB6_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB6), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB6), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTB7,
        GlitchData    => DOUTB7_GlitchData,
        OutSignalName => "DOUTB7",
        OutTemp       => DOUTB7_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB7), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB7), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  VitalPathDelay01Z (
        OutSignal     => DOUTB8,
        GlitchData    => DOUTB8_GlitchData,
        OutSignalName => "DOUTB8",
        OutTemp       => DOUTB8_zd,
        Paths         => (0 => (CLKB_ipd'last_event,
                                VitalExtendToFillDelay(tpd_CLKB_DOUTB8), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_DOUTB8), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );
   
  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_RAM4K9_VITAL of RAM4K9 is
   for VITAL_ACT
   end for;
end CFG_RAM4K9_VITAL;


----- CELL RAM512X18 -----
library IEEE;
library STD;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_timing.all;
use IEEE.VITAL_primitives.all;


use std.textio.all;
use ieee.std_logic_textio.all;

-- entity declaration --
 entity RAM512X18 is
   generic (
      TimingChecksOn  : Boolean := True;
      InstancePath    : String  := "*";
      Xon             : Boolean := False;
      MsgOn           : Boolean := True;
      MEMORYFILE      : String  := "";
      WARNING_MSGS_ON : Boolean := True;

      tipd_RADDR8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RADDR0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR8    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR7    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR6    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR5    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR4    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR3    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR2    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR1    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WADDR0    : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD17      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD16      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD15      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD14      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD13      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD12      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD11      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD10      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD9       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD8       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD7       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD6       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD5       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD4       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD3       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD2       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW1       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW0       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WEN       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WCLK      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REN       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RCLK      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PIPE      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RESET     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      
      tpd_RCLK_RD17  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RCLK_RD16  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD15  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD14  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD13  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD12  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD11  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD10  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD9   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD8   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD7   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD6   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD5   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD4   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD3   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD2   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD1   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD0   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD17 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD16 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD15 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD14 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD13 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD12 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD11 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD10 : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD9  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD8  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD7  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD6  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD5  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD4  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD3  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD2  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD1  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD0  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      
      tsetup_WD17_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD17_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD16_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD16_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD15_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD15_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD14_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD14_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD13_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD13_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD12_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD12_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD11_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD11_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD10_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD10_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WD9_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD9_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD8_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD8_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD7_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD7_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD6_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD6_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD5_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD5_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD4_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD4_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WD0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD17_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD17_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD16_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD16_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD15_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD15_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD14_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD14_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD13_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD13_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD12_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD12_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD11_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD11_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD10_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD10_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WD9_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD9_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD8_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD8_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD7_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD7_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD6_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD6_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD5_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD5_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD4_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD4_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD3_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD3_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD2_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD2_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD1_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD1_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD0_WCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_WD0_WCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_WADDR8_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR8_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR7_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR7_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR6_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR6_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR5_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR5_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR4_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR4_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR3_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR3_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR2_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR2_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR1_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR1_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR0_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_WADDR0_WCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_WADDR8_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;    
      thold_WADDR8_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR7_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR7_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR6_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR6_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR5_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR5_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR4_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR4_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR3_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR3_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR2_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR2_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR1_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR1_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR0_WCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_WADDR0_WCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_WW1_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WW1_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WW0_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WW0_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WEN_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_WEN_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_WW1_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WW1_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WW0_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WW0_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WEN_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WEN_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_RADDR8_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;    
      tsetup_RADDR8_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR7_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR7_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR6_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR6_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR5_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR5_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR4_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR4_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR3_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR3_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR2_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR2_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR1_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR1_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR0_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_RADDR0_RCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_RADDR8_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;    
      thold_RADDR8_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR7_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR7_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR6_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR6_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR5_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR5_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR4_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR4_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR3_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR3_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR2_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR2_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR1_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR1_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR0_RCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_RADDR0_RCLK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_RW1_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_RW1_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_RW0_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_RW0_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_REN_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_REN_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_RW1_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RW1_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RW0_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RW0_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_REN_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_REN_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;      
      tsetup_PIPE_RCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_PIPE_RCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_PIPE_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_PIPE_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tpw_WCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_WCLK_negedge                   : VitalDelayType := 0.000 ns;
      tpw_RCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_RCLK_negedge                   : VitalDelayType := 0.000 ns;
      trecovery_RESET_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      trecovery_RESET_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_RESET_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RESET_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tpw_RESET_negedge                    : VitalDelayType := 0.000 ns
     );

     port (
           RADDR8        : IN STD_ULOGIC ;
           RADDR7        : IN STD_ULOGIC ;
           RADDR6        : IN STD_ULOGIC ;
           RADDR5        : IN STD_ULOGIC ;
           RADDR4        : IN STD_ULOGIC ;
           RADDR3        : IN STD_ULOGIC ;
           RADDR2        : IN STD_ULOGIC ;
           RADDR1        : IN STD_ULOGIC ;  
           RADDR0        : IN STD_ULOGIC ;
           WADDR8        : IN STD_ULOGIC ;
           WADDR7        : IN STD_ULOGIC ;
           WADDR6        : IN STD_ULOGIC ;
           WADDR5        : IN STD_ULOGIC ;
           WADDR4        : IN STD_ULOGIC ;
           WADDR3        : IN STD_ULOGIC ;
           WADDR2        : IN STD_ULOGIC ;
           WADDR1        : IN STD_ULOGIC ;
           WADDR0        : IN STD_ULOGIC ;
           WD17          : IN STD_ULOGIC ;
           WD16          : IN STD_ULOGIC ;
           WD15          : IN STD_ULOGIC ;
           WD14          : IN STD_ULOGIC ;
           WD13          : IN STD_ULOGIC ;
           WD12          : IN STD_ULOGIC ;
           WD11          : IN STD_ULOGIC ;
           WD10          : IN STD_ULOGIC ;
           WD9           : IN STD_ULOGIC ;
           WD8           : IN STD_ULOGIC ;
           WD7           : IN STD_ULOGIC ;
           WD6           : IN STD_ULOGIC ;
           WD5           : IN STD_ULOGIC ;
           WD4           : IN STD_ULOGIC ;
           WD3           : IN STD_ULOGIC ;
           WD2           : IN STD_ULOGIC ;
           WD1           : IN STD_ULOGIC ;
           WD0           : IN STD_ULOGIC ;
           WW1           : IN STD_ULOGIC ;
           WW0           : IN STD_ULOGIC ;
           WEN           : IN STD_ULOGIC ;
           WCLK          : IN STD_ULOGIC ;
           RW1           : IN STD_ULOGIC ;
           RW0           : IN STD_ULOGIC ;
           REN           : IN STD_ULOGIC ;
           RCLK          : IN STD_ULOGIC ;
           PIPE          : IN STD_ULOGIC ;
           RESET         : IN STD_ULOGIC ;
           RD17          : OUT STD_ULOGIC ;
           RD16          : OUT STD_ULOGIC ;
           RD15          : OUT STD_ULOGIC ;
           RD14          : OUT STD_ULOGIC ;
           RD13          : OUT STD_ULOGIC ;
           RD12          : OUT STD_ULOGIC ;
           RD11          : OUT STD_ULOGIC ;
           RD10          : OUT STD_ULOGIC ;
           RD9           : OUT STD_ULOGIC ;
           RD8           : OUT STD_ULOGIC ;
           RD7           : OUT STD_ULOGIC ;
           RD6           : OUT STD_ULOGIC ;
           RD5           : OUT STD_ULOGIC ;
           RD4           : OUT STD_ULOGIC ;
           RD3           : OUT STD_ULOGIC ;
           RD2           : OUT STD_ULOGIC ;
           RD1           : OUT STD_ULOGIC ;
           RD0           : OUT STD_ULOGIC
  );
  attribute VITAL_LEVEL0 of RAM512X18 : entity is TRUE;

end RAM512X18;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM512X18 is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal RADDR8_ipd : std_ulogic := 'X';
  signal RADDR7_ipd : std_ulogic := 'X';
  signal RADDR6_ipd : std_ulogic := 'X';
  signal RADDR5_ipd : std_ulogic := 'X';
  signal RADDR4_ipd : std_ulogic := 'X';
  signal RADDR3_ipd : std_ulogic := 'X';
  signal RADDR2_ipd : std_ulogic := 'X';
  signal RADDR1_ipd : std_ulogic := 'X';
  signal RADDR0_ipd : std_ulogic := 'X';
  signal WADDR8_ipd : std_ulogic := 'X';
  signal WADDR7_ipd : std_ulogic := 'X';
  signal WADDR6_ipd : std_ulogic := 'X';
  signal WADDR5_ipd : std_ulogic := 'X';
  signal WADDR4_ipd : std_ulogic := 'X';
  signal WADDR3_ipd : std_ulogic := 'X';
  signal WADDR2_ipd : std_ulogic := 'X'; 
  signal WADDR1_ipd : std_ulogic := 'X';
  signal WADDR0_ipd : std_ulogic := 'X';
  signal WD17_ipd   : std_ulogic := 'X';
  signal WD16_ipd   : std_ulogic := 'X';
  signal WD15_ipd   : std_ulogic := 'X';
  signal WD14_ipd   : std_ulogic := 'X';
  signal WD13_ipd   : std_ulogic := 'X';
  signal WD12_ipd   : std_ulogic := 'X';
  signal WD11_ipd   : std_ulogic := 'X'; 
  signal WD10_ipd   : std_ulogic := 'X';
  signal WD9_ipd    : std_ulogic := 'X';
  signal WD8_ipd    : std_ulogic := 'X';
  signal WD7_ipd    : std_ulogic := 'X';
  signal WD6_ipd    : std_ulogic := 'X';
  signal WD5_ipd    : std_ulogic := 'X';
  signal WD4_ipd    : std_ulogic := 'X';
  signal WD3_ipd    : std_ulogic := 'X';
  signal WD2_ipd    : std_ulogic := 'X'; 
  signal WD1_ipd    : std_ulogic := 'X';
  signal WD0_ipd    : std_ulogic := 'X';
  signal WW1_ipd    : std_ulogic := 'X';
  signal WW0_ipd    : std_ulogic := 'X';
  signal WEN_ipd    : std_ulogic := 'X'; 
  signal WCLK_ipd   : std_ulogic := 'X';
  signal REN_ipd    : std_ulogic := 'X';
  signal PIPE_ipd   : std_ulogic := 'X';
  signal RESET_ipd  : std_ulogic := 'X';
  signal RW1_ipd    : std_ulogic := 'X'; 
  signal RW0_ipd    : std_ulogic := 'X';
  signal RCLK_ipd   : std_ulogic := 'X'; 
  
  signal INIT_MEM   : std_logic  := '0';       

  type MEMORY_512_9 is array ( 0 to 511, 8 downto 0 ) of std_ulogic; -- memory array with pre-load capability

  constant TC2CWRH   : time       := 1.043 ns;
  constant TC2CRWH   : time       := 0.871 ns;

  -- function to check if write and read operations are accessing the same memory location

  function same_addr(
    waddr, raddr : integer;
    ww, rw       : integer ) return boolean is
    variable result           : boolean;
    variable wr_addr, rd_addr : integer;
  begin
    result := false;

    if ( ww > rw ) then
      rd_addr := ( raddr / (2 ** (ww-rw)) );
      wr_addr := waddr;
    elsif ( rw > ww ) then
      rd_addr := raddr;
      wr_addr := ( waddr / (2 ** (rw-ww)) );
    else
      rd_addr := raddr;
      wr_addr := waddr;
    end if;

    if ( wr_addr = rd_addr ) then
      result := true;
    end if;

    return result;
  end function same_addr;

  -- function to drive read data bus to "x" depending on width configuration

  function drive_rd_x(
    waddr, raddr : integer;
    ww, rw       : integer;
    rd_data      : std_logic_vector (17 downto 0) ) return std_logic_vector is

    variable data_x : std_logic_vector (17 downto 0);
    variable index  : integer;

  begin
    data_x := rd_data;

    case (rw) is
      when 1 =>
              data_x ( 8 downto 0 ) := ( others => 'X' );
      when 2 =>
            if ( ww = 1 ) then
              index := ( waddr mod 2 ) * 9;
              for i in index to index+8 loop
                data_x ( i ) := 'X';
              end loop;
            else
              data_x ( 17 downto 0 ) := ( others => 'X' );
            end if;
      when others =>
            if ( WARNING_MSGS_ON ) then
              assert false
                report "Illegal Read port width configuration"
                severity warning;
            end if;
     end case;

    return data_x;

  end function drive_rd_x;


begin  --  VITAL_ACT

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WireDelay: block

  begin  --  block WireDelay
    VitalWireDelay (RADDR8_ipd, RADDR8, VitalExtendToFillDelay(tipd_RADDR8));
    VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
    VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
    VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
    VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
    VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
    VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
    VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
    VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
    VitalWireDelay (WADDR8_ipd, WADDR8, VitalExtendToFillDelay(tipd_WADDR8));
    VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
    VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
    VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
    VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
    VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
    VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
    VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
    VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
    VitalWireDelay (WD0_ipd,    WD0,    VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (WD1_ipd,    WD1,    VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD2_ipd,    WD2,    VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD3_ipd,    WD3,    VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD4_ipd,    WD4,    VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD5_ipd,    WD5,    VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD6_ipd,    WD6,    VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD7_ipd,    WD7,    VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD8_ipd,    WD8,    VitalExtendToFillDelay(tipd_WD8));
    VitalWireDelay (WD9_ipd,    WD9,    VitalExtendToFillDelay(tipd_WD9));
    VitalWireDelay (WD10_ipd,   WD10,   VitalExtendToFillDelay(tipd_WD10));
    VitalWireDelay (WD11_ipd,   WD11,   VitalExtendToFillDelay(tipd_WD11));
    VitalWireDelay (WD12_ipd,   WD12,   VitalExtendToFillDelay(tipd_WD12));
    VitalWireDelay (WD13_ipd,   WD13,   VitalExtendToFillDelay(tipd_WD13));
    VitalWireDelay (WD14_ipd,   WD14,   VitalExtendToFillDelay(tipd_WD14));
    VitalWireDelay (WD15_ipd,   WD15,   VitalExtendToFillDelay(tipd_WD15));
    VitalWireDelay (WD16_ipd,   WD16,   VitalExtendToFillDelay(tipd_WD16));
    VitalWireDelay (WD17_ipd,   WD17,   VitalExtendToFillDelay(tipd_WD17));
    VitalWireDelay (WW1_ipd,    WW1,    VitalExtendToFillDelay(tipd_WW1));
    VitalWireDelay (WW0_ipd,    WW0,    VitalExtendToFillDelay(tipd_WW0));
    VitalWireDelay (WEN_ipd,    WEN,    VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd,   WCLK,   VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RESET_ipd,  RESET,  VitalExtendToFillDelay(tipd_RESET));
    VitalWireDelay (PIPE_ipd,   PIPE,   VitalExtendToFillDelay(tipd_PIPE));
    VitalWireDelay (REN_ipd,    REN,    VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RW1_ipd,    RW1,    VitalExtendToFillDelay(tipd_RW1));
    VitalWireDelay (RW0_ipd,    RW0,    VitalExtendToFillDelay(tipd_RW0));
    VitalWireDelay (RCLK_ipd,   RCLK,   VitalExtendToFillDelay(tipd_RCLK));

  end block WireDelay;

  -- INITIALIZE MEMORY --

  process
  begin
    INIT_MEM <= '1';
    wait;
  end process;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################
  VITALBehavior : process (RCLK_ipd, REN_ipd, PIPE_ipd, RW1_ipd, RW0_ipd, 
                           WEN_ipd, WCLK_ipd, RESET_ipd, WW1_ipd, WW0_ipd,
                           RADDR8_ipd, RADDR7_ipd, RADDR6_ipd, RADDR5_ipd, 
                           RADDR4_ipd, RADDR3_ipd, RADDR2_ipd, RADDR1_ipd,
                           RADDR0_ipd, WADDR8_ipd, WADDR7_ipd, WADDR6_ipd,
                           WADDR5_ipd, WADDR4_ipd, WADDR3_ipd, WADDR2_ipd,
                           WADDR1_ipd, WADDR0_ipd, WD17_ipd, WD16_ipd,
                           WD15_ipd, WD14_ipd, WD13_ipd, WD12_ipd, WD11_ipd,
                           WD10_ipd, WD9_ipd, WD8_ipd, WD7_ipd, WD6_ipd,
                           WD5_ipd, WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd,
                           WD0_ipd, INIT_MEM)


     -- some internal veriable declaration
     variable RADDR  : integer := 0;
     variable WADDR  : integer := 0;
     variable rwidth : integer := 0;
     variable wwidth : integer := 0;

     variable RADDR_VALID : integer := 1;
     variable WADDR_VALID : integer := 1;

     variable MEM_512_9 : MEMORY_512_9;

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);

     variable i              : integer := 0;
     file     memfile        : text;
     variable status         : file_open_status;
     variable msgs_checked   : Boolean := False;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-511, -511, 0, 1, -511, -511, 0, 1, -511);

     --  Read Timing Check Results
     variable Tviol_WD17_WCLK_posedge : X01 := '0';
     variable TmDt_WD17_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD16_WCLK_posedge : X01 := '0';
     variable TmDt_WD16_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD15_WCLK_posedge : X01 := '0';
     variable TmDt_WD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD14_WCLK_posedge : X01 := '0';
     variable TmDt_WD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD13_WCLK_posedge : X01 := '0';
     variable TmDt_WD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD12_WCLK_posedge : X01 := '0';
     variable TmDt_WD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD11_WCLK_posedge : X01 := '0';
     variable TmDt_WD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD10_WCLK_posedge : X01 := '0';
     variable TmDt_WD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD9_WCLK_posedge : X01 := '0';
     variable TmDt_WD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD8_WCLK_posedge : X01 := '0';
     variable TmDt_WD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW1_WCLK_posedge : X01 := '0';
     variable TmDt_WW1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW0_WCLK_posedge : X01 := '0';
     variable TmDt_WW0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR8_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WCLK_posedge : X01 := '0';
     variable TmDt_WADDR0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR8_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR8_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR7_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR6_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_RCLK_posedge : X01 := '0';
     variable TmDt_RADDR0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PIPE_RCLK_posedge : X01 := '0';
     variable TmDt_PIPE_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW1_RCLK_posedge : X01 := '0';
     variable TmDt_RW1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW0_RCLK_posedge : X01 := '0';
     variable TmDt_RW0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
     variable PeriodData_RESET : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET : X01 := '0';
     variable Tviol_RESET_RCLK_posedge : X01 := '0';
     variable Tmkr_RESET_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLK_posedge : X01 := '0';
     variable Tmkr_RESET_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     
   -- functional Results

     variable RD0_zd   : std_ulogic;
     variable RD1_zd   : std_ulogic;
     variable RD2_zd   : std_ulogic;
     variable RD3_zd   : std_ulogic;
     variable RD4_zd   : std_ulogic;
     variable RD5_zd   : std_ulogic;
     variable RD6_zd   : std_ulogic;
     variable RD7_zd   : std_ulogic;
     variable RD8_zd   : std_ulogic;
     variable RD9_zd   : std_ulogic;
     variable RD10_zd  : std_ulogic;
     variable RD11_zd  : std_ulogic;
     variable RD12_zd  : std_ulogic;
     variable RD13_zd  : std_ulogic;
     variable RD14_zd  : std_ulogic;
     variable RD15_zd  : std_ulogic;
     variable RD16_zd  : std_ulogic;
     variable RD17_zd  : std_ulogic;

     variable RD0_stg  : std_ulogic;
     variable RD1_stg  : std_ulogic;
     variable RD2_stg  : std_ulogic;
     variable RD3_stg  : std_ulogic;
     variable RD4_stg  : std_ulogic;
     variable RD5_stg  : std_ulogic;
     variable RD6_stg  : std_ulogic;
     variable RD7_stg  : std_ulogic;
     variable RD8_stg  : std_ulogic;
     variable RD9_stg  : std_ulogic;
     variable RD10_stg : std_ulogic;
     variable RD11_stg : std_ulogic;
     variable RD12_stg : std_ulogic;
     variable RD13_stg : std_ulogic;
     variable RD14_stg : std_ulogic;
     variable RD15_stg : std_ulogic;
     variable RD16_stg : std_ulogic;
     variable RD17_stg : std_ulogic;


   -- Output Glitch Detection Support Variables

     variable RD0_GlitchData  : VitalGlitchDataType;
     variable RD1_GlitchData  : VitalGlitchDataType;
     variable RD2_GlitchData  : VitalGlitchDataType;
     variable RD3_GlitchData  : VitalGlitchDataType;
     variable RD4_GlitchData  : VitalGlitchDataType;
     variable RD5_GlitchData  : VitalGlitchDataType;
     variable RD6_GlitchData  : VitalGlitchDataType;
     variable RD7_GlitchData  : VitalGlitchDataType;
     variable RD8_GlitchData  : VitalGlitchDataType;
     variable RD9_GlitchData  : VitalGlitchDataType;
     variable RD10_GlitchData : VitalGlitchDataType;
     variable RD11_GlitchData : VitalGlitchDataType;
     variable RD12_GlitchData : VitalGlitchDataType;
     variable RD13_GlitchData : VitalGlitchDataType;
     variable RD14_GlitchData : VitalGlitchDataType;
     variable RD15_GlitchData : VitalGlitchDataType;
     variable RD16_GlitchData : VitalGlitchDataType;
     variable RD17_GlitchData : VitalGlitchDataType;

  
     -- last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';

     variable REN_delayed     : std_ulogic := 'X';
     variable WEN_delayed     : std_ulogic := 'X';
     variable RPIPE_delayed   : std_ulogic := 'X';
     variable RESET_delayed   : std_ulogic := 'X';
     variable WD0_delayed     : std_ulogic := 'X';
     variable WD1_delayed     : std_ulogic := 'X';
     variable WD2_delayed     : std_ulogic := 'X';
     variable WD3_delayed     : std_ulogic := 'X';
     variable WD4_delayed     : std_ulogic := 'X';
     variable WD5_delayed     : std_ulogic := 'X';
     variable WD6_delayed     : std_ulogic := 'X';
     variable WD7_delayed     : std_ulogic := 'X';
     variable WD8_delayed     : std_ulogic := 'X';
     variable WD9_delayed     : std_ulogic := 'X';
     variable WD10_delayed    : std_ulogic := 'X';
     variable WD11_delayed    : std_ulogic := 'X';
     variable WD12_delayed    : std_ulogic := 'X';
     variable WD13_delayed    : std_ulogic := 'X';
     variable WD14_delayed    : std_ulogic := 'X';
     variable WD15_delayed    : std_ulogic := 'X';
     variable WD16_delayed    : std_ulogic := 'X';
     variable WD17_delayed    : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR8_delayed  : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR8_delayed  : std_ulogic := 'X';
    
     -- simultaneous write and read logic detection 

     variable WEN_lat         : std_logic;
     variable REN_lat         : std_logic;
     variable WW_INT          : integer := 0;
     variable RW_INT          : integer := 0;
     variable WCLK_re         : Time;
     variable RCLK_re         : Time;
     variable RD_array        : std_logic_vector ( 17 downto 0 );
  
begin -- process VITALBehavior

  if ( msgs_checked = False ) then
    msgs_checked := True;
    if ( WARNING_MSGS_ON = False ) then
      report "RAM512X18 warnings disabled. Set WARNING_MSGS_ON => True to enable."
      severity note;
    end if;
  end if;
  

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'event and INIT_MEM = '1' ) then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while (( i <= 511 ) and ( not endfile(memfile))) loop
        readline(memfile, inline);
        read(inline, indata);
        resdata := indata;
        MEM_512_9(i,8) := resdata(8);
        MEM_512_9(i,7) := resdata(7);
        MEM_512_9(i,6) := resdata(6);
        MEM_512_9(i,5) := resdata(5);
        MEM_512_9(i,4) := resdata(4);
        MEM_512_9(i,3) := resdata(3);
        MEM_512_9(i,2) := resdata(2);
        MEM_512_9(i,1) := resdata(1);
        MEM_512_9(i,0) := resdata(0);
        i := i + 1;
      end loop;
    else
      if ( WARNING_MSGS_ON ) then
        assert ( MEMORYFILE'length = 0 )
          report "Failed to open memory initialization in read mode"
          severity note;
      end if;
    end if;
    file_close(memfile);
  end if;


  if (TimingChecksOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

  -- recovery / removal check for RCLK to RESET signal ;
     VitalRecoveryRemovalCheck  (
         Violation              => Tviol_RESET_RCLK_posedge,
         TimingData             => Tmkr_RESET_RCLK_posedge,
         TestSignal             => RESET_ipd,
         TestSignalName         => "RESET",
         TestDelay              => 0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0 ns,
         Recovery               => trecovery_RESET_RCLK_posedge_posedge,
         Removal                => thold_RESET_RCLK_posedge_posedge,
         ActiveLow              => TRUE,
         CheckEnabled           => (TO_X01(REN_ipd) = '0'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- recovery / removal check for WCLK to RESET signal ; 
     VitalRecoveryRemovalCheck  (
         Violation              => Tviol_RESET_WCLK_posedge,
         TimingData             => Tmkr_RESET_WCLK_posedge,
         TestSignal             => RESET_ipd,
         TestSignalName         => "RESET",
         TestDelay              => 0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0 ns,
         Recovery               => trecovery_RESET_WCLK_posedge_posedge,
         Removal                => thold_RESET_WCLK_posedge_posedge,
         ActiveLow              => TRUE,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- setup / hold REN, PIPE low when RCLK rising
     VitalSetupHoldCheck ( 
         Violation              => Tviol_REN_RCLK_posedge,
         TimingData             => TmDt_REN_RCLK_posedge,
         TestSignal             => REN_ipd, 
         TestSignalName         => "REN",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_REN_RCLK_posedge_posedge,
         SetupLow               => tsetup_REN_RCLK_negedge_posedge,
         HoldHigh               => thold_REN_RCLK_posedge_posedge,
         HoldLow                => thold_REN_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_PIPE_RCLK_posedge,
         TimingData             => TmDt_PIPE_RCLK_posedge,
         TestSignal             => PIPE_ipd,
         TestSignalName         => "PIPE",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_PIPE_RCLK_posedge_posedge,
         SetupLow               => tsetup_PIPE_RCLK_negedge_posedge,
         HoldHigh               => thold_PIPE_RCLK_posedge_posedge,
         HoldLow                => thold_PIPE_RCLK_negedge_posedge,
         CheckEnabled           => ((TO_X01(RESET_ipd) = '1') and (TO_X01(REN_ipd) ='0')),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- setup / hold WEN when WCLK rising
     VitalSetupHoldCheck ( 
         Violation              => Tviol_WEN_WCLK_posedge,
         TimingData             => TmDt_WEN_WCLK_posedge,
         TestSignal             => WEN_ipd,
         TestSignalName         => "WEN",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WEN_WCLK_posedge_posedge,
         SetupLow               => tsetup_WEN_WCLK_negedge_posedge,
         HoldHigh               => thold_WEN_WCLK_posedge_posedge,
         HoldLow                => thold_WEN_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- setup / hold WD0 - 17 when WCLK rising
     VitalSetupHoldCheck ( 
         Violation              => Tviol_WD0_WCLK_posedge,
         TimingData             => TmDt_WD0_WCLK_posedge,
         TestSignal             => WD0_ipd,
         TestSignalName         => "WD0",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD0_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD0_WCLK_negedge_posedge,
         HoldHigh               => thold_WD0_WCLK_posedge_posedge,
         HoldLow                => thold_WD0_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_WD1_WCLK_posedge,
         TimingData             => TmDt_WD1_WCLK_posedge,
         TestSignal             => WD1_ipd,
         TestSignalName         => "WD1",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD1_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD1_WCLK_negedge_posedge,
         HoldHigh               => thold_WD1_WCLK_posedge_posedge,
         HoldLow                => thold_WD1_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     VitalSetupHoldCheck ( 
         Violation              => Tviol_WD2_WCLK_posedge,
         TimingData             => TmDt_WD2_WCLK_posedge,
         TestSignal             => WD2_ipd,
         TestSignalName         => "WD2",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD2_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD2_WCLK_negedge_posedge,
         HoldHigh               => thold_WD2_WCLK_posedge_posedge,
         HoldLow                => thold_WD2_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck ( 
         Violation              => Tviol_WD3_WCLK_posedge,
         TimingData             => TmDt_WD3_WCLK_posedge,
         TestSignal             => WD3_ipd,
         TestSignalName         => "WD3",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD3_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD3_WCLK_negedge_posedge,
         HoldHigh               => thold_WD3_WCLK_posedge_posedge,
         HoldLow                => thold_WD3_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck ( 
         Violation              => Tviol_WD4_WCLK_posedge,
         TimingData             => TmDt_WD4_WCLK_posedge,
         TestSignal             => WD4_ipd,
         TestSignalName         => "WD4",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD4_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD4_WCLK_negedge_posedge,
         HoldHigh               => thold_WD4_WCLK_posedge_posedge,
         HoldLow                => thold_WD4_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck ( 
         Violation              => Tviol_WD5_WCLK_posedge,
         TimingData             => TmDt_WD5_WCLK_posedge,
         TestSignal             => WD5_ipd,
         TestSignalName         => "WD5",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD5_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD5_WCLK_negedge_posedge,
         HoldHigh               => thold_WD5_WCLK_posedge_posedge,
         HoldLow                => thold_WD5_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD6_WCLK_posedge,
         TimingData             => TmDt_WD6_WCLK_posedge,
         TestSignal             => WD6_ipd,
         TestSignalName         => "WD6",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD6_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD6_WCLK_negedge_posedge,
         HoldHigh               => thold_WD6_WCLK_posedge_posedge,
         HoldLow                => thold_WD6_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD7_WCLK_posedge,
         TimingData             => TmDt_WD7_WCLK_posedge,
         TestSignal             => WD7_ipd,
         TestSignalName         => "WD7",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD7_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD7_WCLK_negedge_posedge,
         HoldHigh               => thold_WD7_WCLK_posedge_posedge,
         HoldLow                => thold_WD7_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD8_WCLK_posedge,
         TimingData             => TmDt_WD8_WCLK_posedge,
         TestSignal             => WD8_ipd,
         TestSignalName         => "WD8",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD8_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD8_WCLK_negedge_posedge,
         HoldHigh               => thold_WD8_WCLK_posedge_posedge,
         HoldLow                => thold_WD8_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD9_WCLK_posedge,
         TimingData             => TmDt_WD9_WCLK_posedge,
         TestSignal             => WD9_ipd,
         TestSignalName         => "WD9",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD9_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD9_WCLK_negedge_posedge,
         HoldHigh               => thold_WD9_WCLK_posedge_posedge,
         HoldLow                => thold_WD9_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD10_WCLK_posedge,
         TimingData             => TmDt_WD10_WCLK_posedge,
         TestSignal             => WD10_ipd,
         TestSignalName         => "WD10",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD10_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD10_WCLK_negedge_posedge,
         HoldHigh               => thold_WD10_WCLK_posedge_posedge,
         HoldLow                => thold_WD10_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD11_WCLK_posedge,
         TimingData             => TmDt_WD11_WCLK_posedge,
         TestSignal             => WD11_ipd,
         TestSignalName         => "WD11",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD11_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD11_WCLK_negedge_posedge,
         HoldHigh               => thold_WD11_WCLK_posedge_posedge,
         HoldLow                => thold_WD11_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD12_WCLK_posedge,
         TimingData             => TmDt_WD12_WCLK_posedge,
         TestSignal             => WD12_ipd,
         TestSignalName         => "WD12",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD12_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD12_WCLK_negedge_posedge,
         HoldHigh               => thold_WD12_WCLK_posedge_posedge,
         HoldLow                => thold_WD12_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD13_WCLK_posedge,
         TimingData             => TmDt_WD13_WCLK_posedge,
         TestSignal             => WD13_ipd,
         TestSignalName         => "WD13",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD13_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD13_WCLK_negedge_posedge,
         HoldHigh               => thold_WD13_WCLK_posedge_posedge,
         HoldLow                => thold_WD13_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD14_WCLK_posedge,
         TimingData             => TmDt_WD14_WCLK_posedge,
         TestSignal             => WD14_ipd,
         TestSignalName         => "WD14",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD14_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD14_WCLK_negedge_posedge,
         HoldHigh               => thold_WD14_WCLK_posedge_posedge,
         HoldLow                => thold_WD14_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD15_WCLK_posedge,
         TimingData             => TmDt_WD15_WCLK_posedge,
         TestSignal             => WD15_ipd,
         TestSignalName         => "WD15",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD15_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD15_WCLK_negedge_posedge,
         HoldHigh               => thold_WD15_WCLK_posedge_posedge,
         HoldLow                => thold_WD15_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD16_WCLK_posedge,
         TimingData             => TmDt_WD16_WCLK_posedge,
         TestSignal             => WD16_ipd,
         TestSignalName         => "WD16",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD16_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD16_WCLK_negedge_posedge,
         HoldHigh               => thold_WD16_WCLK_posedge_posedge,
         HoldLow                => thold_WD16_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WD17_WCLK_posedge,
         TimingData             => TmDt_WD17_WCLK_posedge,
         TestSignal             => WD17_ipd,
         TestSignalName         => "WD17",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WD17_WCLK_posedge_posedge,
         SetupLow               => tsetup_WD17_WCLK_negedge_posedge,
         HoldHigh               => thold_WD17_WCLK_posedge_posedge,
         HoldLow                => thold_WD17_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- setup / hold WADDR0 - 8 to rising edge of WCLK

     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR8_WCLK_posedge,
         TimingData             => TmDt_WADDR8_WCLK_posedge,
         TestSignal             => WADDR8_ipd,
         TestSignalName         => "WADDR8",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR8_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR8_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR8_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR8_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR7_WCLK_posedge,
         TimingData             => TmDt_WADDR7_WCLK_posedge,
         TestSignal             => WADDR7_ipd,
         TestSignalName         => "WADDR7",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR7_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR7_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR7_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR7_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR6_WCLK_posedge,
         TimingData             => TmDt_WADDR6_WCLK_posedge,
         TestSignal             => WADDR6_ipd,
         TestSignalName         => "WADDR6",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR6_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR6_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR6_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR6_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR5_WCLK_posedge,
         TimingData             => TmDt_WADDR5_WCLK_posedge,
         TestSignal             => WADDR5_ipd,
         TestSignalName         => "WADDR5",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR5_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR5_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR5_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR5_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR4_WCLK_posedge,
         TimingData             => TmDt_WADDR4_WCLK_posedge,
         TestSignal             => WADDR4_ipd,
         TestSignalName         => "WADDR4",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR4_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR4_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR4_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR4_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR3_WCLK_posedge,
         TimingData             => TmDt_WADDR3_WCLK_posedge,
         TestSignal             => WADDR3_ipd,
         TestSignalName         => "WADDR3",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR3_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR3_WCLK_negedge_posedge,
         HoldHigh               =>  thold_WADDR3_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR3_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR2_WCLK_posedge,
         TimingData             => TmDt_WADDR2_WCLK_posedge,
         TestSignal             => WADDR2_ipd,
         TestSignalName         => "WADDR2",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR2_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR2_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR2_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR2_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR1_WCLK_posedge,
         TimingData             => TmDt_WADDR1_WCLK_posedge,
         TestSignal             => WADDR1_ipd,
         TestSignalName         => "WADDR1",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR1_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR1_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR1_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR1_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WADDR0_WCLK_posedge,
         TimingData             => TmDt_WADDR0_WCLK_posedge,
         TestSignal             => WADDR0_ipd,
         TestSignalName         => "WADDR0",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WADDR0_WCLK_posedge_posedge,
         SetupLow               => tsetup_WADDR0_WCLK_negedge_posedge,
         HoldHigh               => thold_WADDR0_WCLK_posedge_posedge,
         HoldLow                => thold_WADDR0_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WW0_WCLK_posedge,
         TimingData             => TmDt_WW0_WCLK_posedge,
         TestSignal             => WW0_ipd,
         TestSignalName         => "WW0",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WW0_WCLK_posedge_posedge,
         SetupLow               => tsetup_WW0_WCLK_negedge_posedge,
         HoldHigh               => thold_WW0_WCLK_posedge_posedge,
         HoldLow                => thold_WW0_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_WW1_WCLK_posedge,
         TimingData             => TmDt_WW1_WCLK_posedge,
         TestSignal             => WW1_ipd,
         TestSignalName         => "WW1",
         TestDelay              => 0.0 ns,
         RefSignal              => WCLK_ipd,
         RefSignalName          => "WCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_WW1_WCLK_posedge_posedge,
         SetupLow               => tsetup_WW1_WCLK_negedge_posedge,
         HoldHigh               => thold_WW1_WCLK_posedge_posedge,
         HoldLow                => thold_WW1_WCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR0_RCLK_posedge,
         TimingData             => TmDt_RADDR0_RCLK_posedge,
         TestSignal             => RADDR0_ipd,
         TestSignalName         => "RADDR0",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR0_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR0_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR0_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR0_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR1_RCLK_posedge,
         TimingData             => TmDt_RADDR1_RCLK_posedge,
         TestSignal             => RADDR1_ipd,
         TestSignalName         => "RADDR1",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR1_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR1_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR1_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR1_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR2_RCLK_posedge,
         TimingData             => TmDt_RADDR2_RCLK_posedge,
         TestSignal             => RADDR2_ipd,
         TestSignalName         => "RADDR2",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR2_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR2_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR2_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR2_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR3_RCLK_posedge,
         TimingData             => TmDt_RADDR3_RCLK_posedge,
         TestSignal             => RADDR3_ipd,
         TestSignalName         => "RADDR3",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR3_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR3_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR3_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR3_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR4_RCLK_posedge,
         TimingData             => TmDt_RADDR4_RCLK_posedge,
         TestSignal             => RADDR4_ipd,
         TestSignalName         => "RADDR4",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR4_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR4_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR4_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR4_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR5_RCLK_posedge,
         TimingData             => TmDt_RADDR5_RCLK_posedge,
         TestSignal             => RADDR5_ipd,
         TestSignalName         => "RADDR5",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR5_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR5_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR5_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR5_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR6_RCLK_posedge,
         TimingData             => TmDt_RADDR6_RCLK_posedge,
         TestSignal             => RADDR6_ipd,
         TestSignalName         => "RADDR6",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR6_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR6_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR6_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR6_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR7_RCLK_posedge,
         TimingData             => TmDt_RADDR7_RCLK_posedge,
         TestSignal             => RADDR7_ipd,
         TestSignalName         => "RADDR7",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR7_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR7_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR7_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR7_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RADDR8_RCLK_posedge,
         TimingData             => TmDt_RADDR8_RCLK_posedge,
         TestSignal             => RADDR8_ipd,
         TestSignalName         => "RADDR8",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RADDR8_RCLK_posedge_posedge,
         SetupLow               => tsetup_RADDR8_RCLK_negedge_posedge,
         HoldHigh               => thold_RADDR8_RCLK_posedge_posedge,
         HoldLow                => thold_RADDR8_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RW1_RCLK_posedge,
         TimingData             => TmDt_RW1_RCLK_posedge,
         TestSignal             => RW1_ipd,
         TestSignalName         => "RW1",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RW1_RCLK_posedge_posedge,
         SetupLow               => tsetup_RW1_RCLK_negedge_posedge,
         HoldHigh               => thold_RW1_RCLK_posedge_posedge,
         HoldLow                => thold_RW1_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );
         
     VitalSetupHoldCheck (
         Violation              => Tviol_RW0_RCLK_posedge,
         TimingData             => TmDt_RW0_RCLK_posedge,
         TestSignal             => RW0_ipd,
         TestSignalName         => "RW0",
         TestDelay              => 0.0 ns,
         RefSignal              => RCLK_ipd,
         RefSignalName          => "RCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_RW0_RCLK_posedge_posedge,
         SetupLow               => tsetup_RW0_RCLK_negedge_posedge,
         HoldHigh               => thold_RW0_RCLK_posedge_posedge,
         HoldLow                => thold_RW0_RCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  --   Period of RCLK
     VitalPeriodPulseCheck (
         Violation              => Pviol_RCLK,
         PeriodData             => PeriodData_RCLK,
         TestSignal             => RCLK_ipd,
         TestSignalName         => "RCLK",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => tpw_RCLK_posedge,
         PulseWidthLow          => tpw_RCLK_negedge,
         CheckEnabled           => ((TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  --   Period of WCLK
     VitalPeriodPulseCheck ( 
         Violation              => Pviol_WCLK,
         PeriodData             => PeriodData_WCLK,
         TestSignal             => WCLK_ipd,
         TestSignalName         => "WCLK",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => tpw_WCLK_posedge,
         PulseWidthLow          => tpw_WCLK_negedge,
         CheckEnabled           => ((TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  --   Period of RESET
     VitalPeriodPulseCheck ( 
         Violation              => Pviol_RESET,
         PeriodData             => PeriodData_RESET,
         TestSignal             => RESET_ipd,
         TestSignalName         => "RESET",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => 0.0 ns,
         PulseWidthLow          => tpw_RESET_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/RAM512X18",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     end if;
     
   -----------------------------------------------------------
   --    Calculate the WW and RW values
   -----------------------------------------------------------

   if ( WW1_ipd'event or WW0_ipd'event ) then
     if ((TO_X01(WW1_ipd) = '0') and (TO_X01(WW0_ipd) = '1')) then
       wwidth := 9;
       WW_INT := 1;
     elsif ((TO_X01(WW1_ipd) = '1') and (TO_X01(WW0_ipd) = '0')) then
       wwidth := 18;
       WW_INT := 2;
     else
       wwidth := -1;
       WW_INT := -1;
     end if;
   end if;

   if ( RW1_ipd'event or RW0_ipd'event ) then
     if ((TO_X01(RW1_ipd) = '0') and (TO_X01(RW0_ipd) = '1')) then
       rwidth := 9;
       RW_INT := 1;
     elsif ((TO_X01(RW1_ipd) = '1') and (TO_X01(RW0_ipd) = '0')) then
       rwidth := 18;
       RW_INT := 2;
     else
       rwidth := -1;
       RW_INT := -1;
     end if;
   end if;

  -----------------------------------------------------------
  --    Check if address out of range for specified width  --
  -----------------------------------------------------------
  
  if (TO_X01(RESET_ipd) = '1' and TO_X01(WEN_delayed) = '0') then
    if (WCLK_ipd'event and TO_X01(WCLK_ipd) = '1') then

      WCLK_re := now;

      -- Calculate the integer value of WADDR

      WADDR := (INT(WADDR8_ipd)*256) +
               (INT(WADDR7_ipd)*128) + (INT(WADDR6_ipd)*64) +
               (INT(WADDR5_ipd)*32)  + (INT(WADDR4_ipd)*16) +
               (INT(WADDR3_ipd)*8)   + (INT(WADDR2_ipd)*4)  +
               (INT(WADDR1_ipd)*2)   + (INT(WADDR0_ipd)*1);

      if (WADDR < 0) then
        WADDR_VALID := 0;
      else
        WADDR_VALID := 1;
      end if;

      if (wwidth = 9 and WADDR >= 512) then
        WADDR_VALID := 0;
      elsif (wwidth = 18 and WADDR >= 256) then
        WADDR_VALID := 0;
      end if;

      if ( WARNING_MSGS_ON ) then
        assert (wwidth /= 9 or (WADDR < 512 and WADDR >= 0) )
          report "Illegal address on Write Port, should be between 0 & 511."
          severity Warning;

        assert (wwidth /= 18 or (WADDR < 256 and WADDR >= 0) )
          report "Illegal address on Write port, should be between 0 & 255."
          severity Warning;
      end if;

    end if;
  end if;
  
  if (TO_X01(RESET_ipd) = '1' and TO_X01(REN_delayed) = '0') then
    if (RCLK_ipd'event and TO_X01(RCLK_ipd) = '1') then

      RCLK_re := now;

      -- Calculate the integer value of RADDR

      RADDR := (INT(RADDR8_ipd)*256) +
               (INT(RADDR7_ipd)*128) + (INT(RADDR6_ipd)*64) +
               (INT(RADDR5_ipd)*32)  + (INT(RADDR4_ipd)*16) +
               (INT(RADDR3_ipd)*8)   + (INT(RADDR2_ipd)*4)  +
               (INT(RADDR1_ipd)*2)   + (INT(RADDR0_ipd)*1);

      if (RADDR < 0) then
        RADDR_VALID := 0;
      else
        RADDR_VALID := 1;
      end if;

      if (rwidth = 9 and RADDR >= 512) then
        RADDR_VALID := 0;
      elsif (rwidth = 18 and RADDR >= 256) then
        RADDR_VALID := 0;
      end if;

      if ( WARNING_MSGS_ON ) then
        assert (rwidth /= 9 or (RADDR < 512 and RADDR >= 0) )
          report "Illegal address on Read Port, should be between 0 & 511."
          severity Warning;

        assert (rwidth /= 18 or (RADDR < 256 and RADDR >= 0) )
          report "Illegal address on Read port, should be between 0 & 255."
          severity Warning;
      end if;

    end if;
  end if;

  -----------------------------------------------------------
  --  RAM RESET
  -----------------------------------------------------------

  if (RESET_ipd'event and TO_X01(RESET_ipd) = '0') then
    case (rwidth) is
      when 9  =>
              RD0_zd := '0';
              RD1_zd := '0';
              RD2_zd := '0';
              RD3_zd := '0';
              RD4_zd := '0';
              RD5_zd := '0';
              RD6_zd := '0';
              RD7_zd := '0';
              RD8_zd := '0';
      when 18 =>
              RD0_zd := '0';
              RD1_zd := '0';
              RD2_zd := '0';
              RD3_zd := '0';
              RD4_zd := '0';
              RD5_zd := '0';
              RD6_zd := '0';
              RD7_zd := '0';
              RD8_zd := '0';
              RD9_zd := '0';
              RD10_zd := '0';
              RD11_zd := '0';
              RD12_zd := '0';
              RD13_zd := '0';
              RD14_zd := '0';
              RD15_zd := '0';
              RD16_zd := '0';
              RD17_zd := '0';
      when others =>
             -- if ( WARNING_MSGS_ON ) then
              --  assert false
              --    report "Illegal Read port width configuration"
              --    severity Warning;
             -- end if;
    end case;

    if (TO_X01(PIPE_ipd) = '1') then
      case (rwidth) is
        when 9  =>
              RD0_stg := '0';
              RD1_stg := '0';
              RD2_stg := '0';
              RD3_stg := '0';
              RD4_stg := '0';
              RD5_stg := '0';
              RD6_stg := '0';
              RD7_stg := '0';
              RD8_stg := '0';
        when 18 =>
              RD0_stg := '0';
              RD1_stg := '0';
              RD2_stg := '0';
              RD3_stg := '0';
              RD4_stg := '0';
              RD5_stg := '0';
              RD6_stg := '0';
              RD7_stg := '0';
              RD8_stg := '0';
              RD9_stg := '0';
              RD10_stg := '0';
              RD11_stg := '0';
              RD12_stg := '0';
              RD13_stg := '0';
              RD14_stg := '0';
              RD15_stg := '0';
              RD16_stg := '0';
              RD17_stg := '0';
        when others =>
             -- if ( WARNING_MSGS_ON ) then
             --   assert false
             --     report "Illegal Read port width configuration"
             --     severity Warning;
             -- end if;
      end case;
    end if;
  end if; 

  --------------------------------------------------------------------
  --          RAM256X18 READ SECTION                                --
  --------------------------------------------------------------------

  if (TO_X01(RCLK_ipd) = 'X') then
    if ((TO_X01(REN_ipd) ='0') and (TO_X01(RESET_ipd) = '1')) then
      if (TO_X01(RCLK_previous) /= 'X') then
        if ( WARNING_MSGS_ON ) then
          assert false
            report "RCLK unknown"
            severity Warning;
        end if;
        RD0_zd   := 'X';
        RD1_zd   := 'X';
        RD2_zd   := 'X';
        RD3_zd   := 'X';
        RD4_zd   := 'X';
        RD5_zd   := 'X';
        RD6_zd   := 'X';
        RD7_zd   := 'X';
        RD8_zd   := 'X';
        RD9_zd   := 'X';
        RD10_zd  := 'X';
        RD11_zd  := 'X';
        RD12_zd  := 'X';
        RD13_zd  := 'X';
        RD14_zd  := 'X';
        RD15_zd  := 'X';
        RD16_zd  := 'X';
        RD17_zd  := 'X';
      end if;
    end if;
  elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1') and (TO_X01(RESET_delayed) = '1')) then

      REN_lat := REN_ipd;

      --clocking the pipelined data to read data bus

      if (TO_X01(PIPE_ipd) = '1') then
        case (rwidth) is
          when 9  =>
              RD0_zd := RD0_stg;
              RD1_zd := RD1_stg;
              RD2_zd := RD2_stg;
              RD3_zd := RD3_stg;
              RD4_zd := RD4_stg;
              RD5_zd := RD5_stg;
              RD6_zd := RD6_stg;
              RD7_zd := RD7_stg;
              RD8_zd := RD8_stg;
          when 18 =>
              RD0_zd  := RD0_stg;
              RD1_zd  := RD1_stg;
              RD2_zd  := RD2_stg;
              RD3_zd  := RD3_stg;
              RD4_zd  := RD4_stg;
              RD5_zd  := RD5_stg;
              RD6_zd  := RD6_stg;
              RD7_zd  := RD7_stg;
              RD8_zd  := RD8_stg;
              RD9_zd  := RD9_stg;
              RD10_zd := RD10_stg;
              RD11_zd := RD11_stg;
              RD12_zd := RD12_stg;
              RD13_zd := RD13_stg;
              RD14_zd := RD14_stg;
              RD15_zd := RD15_stg;
              RD16_zd := RD16_stg;
              RD17_zd := RD17_stg;
          when others =>
              if ( WARNING_MSGS_ON ) then
                assert false
                  report ": Illegal Read port width configuration"
                  severity Warning;
              end if;
        end case;
      elsif (TO_X01(PIPE_ipd) = 'X') then
        if ( WARNING_MSGS_ON ) then
          assert false
            report "PIPE signal unknown."
            severity Warning;
        end if;
        RD0_zd  := 'X';
        RD1_zd  := 'X';
        RD2_zd  := 'X';
        RD3_zd  := 'X';
        RD4_zd  := 'X';
        RD5_zd  := 'X';
        RD6_zd  := 'X';
        RD7_zd  := 'X';
        RD8_zd  := 'X';
        RD9_zd  := 'X';
        RD10_zd := 'X';
        RD11_zd := 'X';
        RD12_zd := 'X';
        RD13_zd := 'X';
        RD14_zd := 'X';
        RD15_zd := 'X';
        RD16_zd := 'X';
        RD17_zd := 'X';
      end if;

    if (TO_X01(REN_ipd) ='0') and (RADDR_VALID = 1) then


      if (TO_X01(PIPE_ipd) = '0') then
        case (rwidth) is
          when 9  =>
                RD0_zd := MEM_512_9( (RADDR), 0 );
                RD1_zd := MEM_512_9( (RADDR), 1 );
                RD2_zd := MEM_512_9( (RADDR), 2 );
                RD3_zd := MEM_512_9( (RADDR), 3 );
                RD4_zd := MEM_512_9( (RADDR), 4 );
                RD5_zd := MEM_512_9( (RADDR), 5 );
                RD6_zd := MEM_512_9( (RADDR), 6 );
                RD7_zd := MEM_512_9( (RADDR), 7 );
                RD8_zd := MEM_512_9( (RADDR), 8 );

          when 18 =>
                RD0_zd  := MEM_512_9( (RADDR * 2), 0 );
                RD1_zd  := MEM_512_9( (RADDR * 2), 1 );
                RD2_zd  := MEM_512_9( (RADDR * 2), 2 );
                RD3_zd  := MEM_512_9( (RADDR * 2), 3 );
                RD4_zd  := MEM_512_9( (RADDR * 2), 4 );
                RD5_zd  := MEM_512_9( (RADDR * 2), 5 );
                RD6_zd  := MEM_512_9( (RADDR * 2), 6 );
                RD7_zd  := MEM_512_9( (RADDR * 2), 7 );
                RD8_zd  := MEM_512_9( (RADDR * 2), 8 );
                RD9_zd  := MEM_512_9( (RADDR * 2 + 1), 0 );
                RD10_zd := MEM_512_9( (RADDR * 2 + 1), 1 );
                RD11_zd := MEM_512_9( (RADDR * 2 + 1), 2 );
                RD12_zd := MEM_512_9( (RADDR * 2 + 1), 3 );
                RD13_zd := MEM_512_9( (RADDR * 2 + 1), 4 );
                RD14_zd := MEM_512_9( (RADDR * 2 + 1), 5 );
                RD15_zd := MEM_512_9( (RADDR * 2 + 1), 6 );
                RD16_zd := MEM_512_9( (RADDR * 2 + 1), 7 );
                RD17_zd := MEM_512_9( (RADDR * 2 + 1), 8 );

          when others =>
                if ( WARNING_MSGS_ON ) then
                  assert false
                    report "Illegal Read port width configuration"
                    severity Warning;
                end if;
        end case;

        -- Check for Write and Read to the same address, write is not affected
        if ( (WEN_lat = '0') and same_addr(WADDR, RADDR, WW_INT, RW_INT) and
                                                ((WCLK_re + TC2CWRH) > RCLK_re) ) then
          assert false
          report " Write and Read to same address at same time.  RD is unpredictable, driving RD to X "
          severity warning;

          RD_array := ( RD17_zd & RD16_zd & RD15_zd & RD14_zd & RD13_zd & RD12_zd &
                        RD11_zd & RD10_zd & RD9_zd & RD8_zd & RD7_zd & RD6_zd &
                        RD5_zd & RD4_zd & RD3_zd & RD2_zd & RD1_zd & RD0_zd );

          RD_array := drive_rd_x ( WADDR, RADDR, WW_INT, RW_INT, RD_array );
          RD17_zd  := RD_array (17);
          RD16_zd  := RD_array (16);
          RD15_zd  := RD_array (15);
          RD14_zd  := RD_array (14);
          RD13_zd  := RD_array (13);
          RD12_zd  := RD_array (12);
          RD11_zd  := RD_array (11);
          RD10_zd  := RD_array (10);
          RD9_zd   := RD_array ( 9);
          RD8_zd   := RD_array ( 8);
          RD7_zd   := RD_array ( 7);
          RD6_zd   := RD_array ( 6);
          RD5_zd   := RD_array ( 5);
          RD4_zd   := RD_array ( 4);
          RD3_zd   := RD_array ( 3);
          RD2_zd   := RD_array ( 2);
          RD1_zd   := RD_array ( 1);
          RD0_zd   := RD_array ( 0);
        end if;

      elsif (TO_X01(PIPE_ipd) = '1') then
        case (rwidth) is
          when 9  =>
                RD0_stg := MEM_512_9( (RADDR), 0 );
                RD1_stg := MEM_512_9( (RADDR), 1 );
                RD2_stg := MEM_512_9( (RADDR), 2 );
                RD3_stg := MEM_512_9( (RADDR), 3 );
                RD4_stg := MEM_512_9( (RADDR), 4 );
                RD5_stg := MEM_512_9( (RADDR), 5 );
                RD6_stg := MEM_512_9( (RADDR), 6 );
                RD7_stg := MEM_512_9( (RADDR), 7 );
                RD8_stg := MEM_512_9( (RADDR), 8 );

          when 18 =>
                RD0_stg  := MEM_512_9( (RADDR * 2), 0 );
                RD1_stg  := MEM_512_9( (RADDR * 2), 1 );
                RD2_stg  := MEM_512_9( (RADDR * 2), 2 );
                RD3_stg  := MEM_512_9( (RADDR * 2), 3 );
                RD4_stg  := MEM_512_9( (RADDR * 2), 4 );
                RD5_stg  := MEM_512_9( (RADDR * 2), 5 );
                RD6_stg  := MEM_512_9( (RADDR * 2), 6 );
                RD7_stg  := MEM_512_9( (RADDR * 2), 7 );
                RD8_stg  := MEM_512_9( (RADDR * 2), 8 );
                RD9_stg  := MEM_512_9( (RADDR * 2 + 1), 0 );
                RD10_stg := MEM_512_9( (RADDR * 2 + 1), 1 );
                RD11_stg := MEM_512_9( (RADDR * 2 + 1), 2 );
                RD12_stg := MEM_512_9( (RADDR * 2 + 1), 3 );
                RD13_stg := MEM_512_9( (RADDR * 2 + 1), 4 );
                RD14_stg := MEM_512_9( (RADDR * 2 + 1), 5 );
                RD15_stg := MEM_512_9( (RADDR * 2 + 1), 6 );
                RD16_stg := MEM_512_9( (RADDR * 2 + 1), 7 );
                RD17_stg := MEM_512_9( (RADDR * 2 + 1), 8 );
          when others =>
              if ( WARNING_MSGS_ON ) then
                assert false
                  report ": Illegal Read port width configuration"
                  severity Warning;
              end if;
        end case;

        -- Check for Write and Read to the same address, write is not affected
        if ( (WEN_lat = '0') and same_addr(WADDR, RADDR, WW_INT, RW_INT) and
                                                ((WCLK_re + TC2CWRH) > RCLK_re) ) then

          assert false
          report " Write and Read to same address at same time.  RD is unpredictable, driving RD to X "
          severity warning;

          RD_array := ( RD17_stg & RD16_stg & RD15_stg & RD14_stg & RD13_stg & RD12_stg &
                        RD11_stg & RD10_stg & RD9_stg & RD8_stg & RD7_stg & RD6_stg &
                        RD5_stg & RD4_stg & RD3_stg & RD2_stg & RD1_stg & RD0_stg );
  
          RD_array := drive_rd_x ( WADDR, RADDR, WW_INT, RW_INT, RD_array );
          RD17_stg := RD_array (17);
          RD16_stg := RD_array (16);
          RD15_stg := RD_array (15);
          RD14_stg := RD_array (14);
          RD13_stg := RD_array (13);
          RD12_stg := RD_array (12);
          RD11_stg := RD_array (11);
          RD10_stg := RD_array (10);
          RD9_stg  := RD_array ( 9);
          RD8_stg  := RD_array ( 8);
          RD7_stg  := RD_array ( 7);
          RD6_stg  := RD_array ( 6);
          RD5_stg  := RD_array ( 5);
          RD4_stg  := RD_array ( 4);
          RD3_stg  := RD_array ( 3);
          RD2_stg  := RD_array ( 2);
          RD1_stg  := RD_array ( 1);
          RD0_stg  := RD_array ( 0);
        end if;

      else
        if ( WARNING_MSGS_ON ) then
          assert false
            report "PIPE signal unknown."
            severity Warning;
        end if;
        RD0_zd  := 'X';
        RD1_zd  := 'X';
        RD2_zd  := 'X';
        RD3_zd  := 'X';
        RD4_zd  := 'X';
        RD5_zd  := 'X';
        RD6_zd  := 'X';
        RD7_zd  := 'X';
        RD8_zd  := 'X';
        RD9_zd  := 'X';
        RD10_zd := 'X';
        RD11_zd := 'X';
        RD12_zd := 'X';
        RD13_zd := 'X';
        RD14_zd := 'X';
        RD15_zd := 'X';
        RD16_zd := 'X';
        RD17_zd := 'X';
      end if;
    elsif (TO_X01(REN_ipd) = '0') and (RADDR_VALID = 0) then
      if ( WARNING_MSGS_ON ) then
        assert false
          report "Illegal Read Address, Read Not Initiated."
          severity Warning;
      end if;
    elsif (TO_X01(REN_ipd) /= '1') then
      if ( WARNING_MSGS_ON ) then
        assert false
          report "REN unknown. "
          severity Warning;
      end if;
    end if;
  end if;

  ------------------------------------------------------------
  -- # Write Functional Section                             --
  ------------------------------------------------------------

  if (TO_X01(WCLK_ipd) = 'X') then
    if ((TO_X01(RESET_ipd) = '1') and (TO_X01(WEN_ipd) = '0')) then 
      if (TO_X01(WCLK_previous) /= 'X') then
        if ( WARNING_MSGS_ON ) then
          assert false
            report "WCLK unknown"
            severity Warning;
        end if;
      end if;
    end if;
  elsif (WCLK_ipd'event and TO_X01(WCLK_ipd) = '1') and (TO_X01(RESET_delayed) = '1') then

    WEN_lat := WEN_ipd;

    if (TO_X01(WEN_ipd) = '0') and (WADDR_VALID = 1) then

      -- Check for Write and Read to the same address, write is not affected
      if ( (REN_lat = '0') and same_addr(WADDR, RADDR, WW_INT, RW_INT) and
                                           ((RCLK_re + TC2CRWH) > WCLK_re) ) then
        assert false
        report " Read and Write to same address at same time.  RD is unpredictable, driving RD to X "
        severity warning;

        if (TO_X01(PIPE_ipd) = '1') then --pipelining on
          RD_array := ( RD17_stg & RD16_stg & RD15_stg & RD14_stg & RD13_stg & RD12_stg &
                        RD11_stg & RD10_stg & RD9_stg & RD8_stg & RD7_stg & RD6_stg &
                        RD5_stg & RD4_stg & RD3_stg & RD2_stg & RD1_stg & RD0_stg );

          -- function call to determine conflicting read data bits based on address and width configuration
          RD_array := drive_rd_x ( WADDR, RADDR, WW_INT, RW_INT, RD_array );

          RD17_stg := RD_array (17);
          RD16_stg := RD_array (16);
          RD15_stg := RD_array (15);
          RD14_stg := RD_array (14);
          RD13_stg := RD_array (13);
          RD12_stg := RD_array (12);
          RD11_stg := RD_array (11);
          RD10_stg := RD_array (10);
          RD9_stg  := RD_array ( 9);
          RD8_stg  := RD_array ( 8);
          RD7_stg  := RD_array ( 7);
          RD6_stg  := RD_array ( 6);
          RD5_stg  := RD_array ( 5);
          RD4_stg  := RD_array ( 4);
          RD3_stg  := RD_array ( 3);
          RD2_stg  := RD_array ( 2);
          RD1_stg  := RD_array ( 1);
          RD0_stg  := RD_array ( 0);
        elsif (TO_X01(PIPE_ipd) = '0') then --pipelining off
          RD_array := ( RD17_zd & RD16_zd & RD15_zd & RD14_zd & RD13_zd & RD12_zd &
                        RD11_zd & RD10_zd & RD9_zd & RD8_zd & RD7_zd & RD6_zd &
                        RD5_zd & RD4_zd & RD3_zd & RD2_zd & RD1_zd & RD0_zd );

          -- function call to determine conflicting read data bits based on address and width configuration
          RD_array := drive_rd_x ( WADDR, RADDR, WW_INT, RW_INT, RD_array );

          RD17_zd  := RD_array (17);
          RD16_zd  := RD_array (16);
          RD15_zd  := RD_array (15);
          RD14_zd  := RD_array (14);
          RD13_zd  := RD_array (13);
          RD12_zd  := RD_array (12);
          RD11_zd  := RD_array (11);
          RD10_zd  := RD_array (10);
          RD9_zd   := RD_array ( 9);
          RD8_zd   := RD_array ( 8);
          RD7_zd   := RD_array ( 7);
          RD6_zd   := RD_array ( 6);
          RD5_zd   := RD_array ( 5);
          RD4_zd   := RD_array ( 4);
          RD3_zd   := RD_array ( 3);
          RD2_zd   := RD_array ( 2);
          RD1_zd   := RD_array ( 1);
          RD0_zd   := RD_array ( 0);
        end if;
      end if;

      -- write data update to memory array
      case(wwidth) is
        when 9 =>
                   MEM_512_9( (WADDR), 0 ) := WD0_delayed;
                   MEM_512_9( (WADDR), 1 ) := WD1_delayed;
                   MEM_512_9( (WADDR), 2 ) := WD2_delayed;
                   MEM_512_9( (WADDR), 3 ) := WD3_delayed;
                   MEM_512_9( (WADDR), 4 ) := WD4_delayed;
                   MEM_512_9( (WADDR), 5 ) := WD5_delayed;
                   MEM_512_9( (WADDR), 6 ) := WD6_delayed;
                   MEM_512_9( (WADDR), 7 ) := WD7_delayed;
                   MEM_512_9( (WADDR), 8 ) := WD8_delayed;
        when 18 =>
                   MEM_512_9( (WADDR * 2), 0 ) := WD0_delayed;
                   MEM_512_9( (WADDR * 2), 1 ) := WD1_delayed;
                   MEM_512_9( (WADDR * 2), 2 ) := WD2_delayed;
                   MEM_512_9( (WADDR * 2), 3 ) := WD3_delayed;
                   MEM_512_9( (WADDR * 2), 4 ) := WD4_delayed;
                   MEM_512_9( (WADDR * 2), 5 ) := WD5_delayed;
                   MEM_512_9( (WADDR * 2), 6 ) := WD6_delayed;
                   MEM_512_9( (WADDR * 2), 7 ) := WD7_delayed;
                   MEM_512_9( (WADDR * 2), 8 ) := WD8_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 0 ) := WD9_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 1 ) := WD10_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 2 ) := WD11_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 3 ) := WD12_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 4 ) := WD13_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 5 ) := WD14_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 6 ) := WD15_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 7 ) := WD16_delayed;
                   MEM_512_9( (WADDR * 2 + 1), 8 ) := WD17_delayed;
        when others =>
                   if ( WARNING_MSGS_ON ) then
                     assert false
                       report "Illegal Write port width configuration"
                       severity Warning;
                   end if;
      end case;
    elsif (TO_X01(WEN_ipd) = '0') and (WADDR_VALID = 0) then
      if ( WARNING_MSGS_ON ) then
        assert false
          report "Illegal Write Address, Write Not Initiated."
          severity Warning;
      end if;
    elsif (TO_X01(WEN_ipd) /= '1') then
      if ( WARNING_MSGS_ON ) then
        assert false
          report "WEN unknown, no data was written into RAM"
          severity Warning;
      end if;
    end if;

  end if;
 
  --------------------------------------------------------------------
  --          Other stuff                                           --
  --------------------------------------------------------------------
 
  if (WCLK_ipd'event) then
     WCLK_previous := WCLK_ipd;
  end if;

  if (RCLK_ipd'event) then
      RCLK_previous := RCLK_ipd;
  end if;
 
                    
  WADDR8_delayed := WADDR8_ipd;
  WADDR7_delayed := WADDR7_ipd;
  WADDR6_delayed := WADDR6_ipd;
  WADDR5_delayed := WADDR5_ipd;
  WADDR4_delayed := WADDR4_ipd;
  WADDR3_delayed := WADDR3_ipd;
  WADDR2_delayed := WADDR2_ipd;
  WADDR1_delayed := WADDR1_ipd;
  WADDR0_delayed := WADDR0_ipd;

  RADDR8_delayed := RADDR8_ipd;
  RADDR7_delayed := RADDR7_ipd;
  RADDR6_delayed := RADDR6_ipd;
  RADDR5_delayed := RADDR5_ipd;
  RADDR4_delayed := RADDR4_ipd;
  RADDR3_delayed := RADDR3_ipd;
  RADDR2_delayed := RADDR2_ipd;
  RADDR1_delayed := RADDR1_ipd;
  RADDR0_delayed := RADDR0_ipd;

  WD17_delayed  := WD17_ipd;
  WD16_delayed  := WD16_ipd;
  WD15_delayed  := WD15_ipd;
  WD14_delayed  := WD14_ipd;
  WD13_delayed  := WD13_ipd;
  WD12_delayed  := WD12_ipd;
  WD11_delayed  := WD11_ipd;
  WD10_delayed  := WD10_ipd;
  WD9_delayed   := WD9_ipd;
  WD8_delayed   := WD8_ipd;
  WD7_delayed   := WD7_ipd;
  WD6_delayed   := WD6_ipd;
  WD5_delayed   := WD5_ipd;
  WD4_delayed   := WD4_ipd;
  WD3_delayed   := WD3_ipd;
  WD2_delayed   := WD2_ipd;
  WD1_delayed   := WD1_ipd;
  WD0_delayed   := WD0_ipd;

  WEN_delayed   := WEN_ipd;
  REN_delayed   := REN_ipd;
  RESET_delayed := RESET_ipd;   
  
  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

    VitalPathDelay01Z (
        OutSignal     => RD17,
        GlitchData    => RD17_GlitchData,
        OutSignalName => "RD17",
        OutTemp       => RD17_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD17), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD17), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD16,
        GlitchData    => RD16_GlitchData,
        OutSignalName => "RD16",
        OutTemp       => RD16_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD16), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD16), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD15,
        GlitchData    => RD15_GlitchData,
        OutSignalName => "RD15",
        OutTemp       => RD15_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD15), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD15), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD14,
        GlitchData    => RD14_GlitchData,
        OutSignalName => "RD14",
        OutTemp       => RD14_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD14), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD14), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD13,
        GlitchData    => RD13_GlitchData,
        OutSignalName => "RD13",
        OutTemp       => RD13_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD13), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD13), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD12,
        GlitchData    => RD12_GlitchData,
        OutSignalName => "RD12",
        OutTemp       => RD12_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD12), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD12), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD11,
        GlitchData    => RD11_GlitchData,
        OutSignalName => "RD11",
        OutTemp       => RD11_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD11), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD11), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD10,
        GlitchData    => RD10_GlitchData,
        OutSignalName => "RD10",
        OutTemp       => RD10_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD10), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD10), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD9,
        GlitchData    => RD9_GlitchData,
        OutSignalName => "RD9",
        OutTemp       => RD9_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD9), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD9), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD8,
        GlitchData    => RD8_GlitchData,
        OutSignalName => "RD8",
        OutTemp       => RD8_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD8), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD8), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD7,
        GlitchData    => RD7_GlitchData,
        OutSignalName => "RD7",
        OutTemp       => RD7_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD7), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD6,
        GlitchData    => RD6_GlitchData,
        OutSignalName => "RD6",
        OutTemp       => RD6_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD6), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD5,
        GlitchData    => RD5_GlitchData,
        OutSignalName => "RD5",
        OutTemp       => RD5_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD5), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD4,
        GlitchData    => RD4_GlitchData,
        OutSignalName => "RD4",
        OutTemp       => RD4_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD4), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD3,
        GlitchData    => RD3_GlitchData,
        OutSignalName => "RD3",
        OutTemp       => RD3_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD3), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD2,
        GlitchData    => RD2_GlitchData,
        OutSignalName => "RD2",
        OutTemp       => RD2_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD2), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD1,
        GlitchData    => RD1_GlitchData,
        OutSignalName => "RD1",
        OutTemp       => RD1_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD1), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

    VitalPathDelay01Z (
        OutSignal     => RD0,
        GlitchData    => RD0_GlitchData,
        OutSignalName => "RD0",
        OutTemp       => RD0_zd,
        Paths         => (0 => (RCLK_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE),
                          1 => (RESET_ipd'last_event,
                                VitalExtendToFillDelay(tpd_RESET_RD0), TRUE)
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );


  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_RAM512X18_VITAL of RAM512X18 is
   for VITAL_ACT
   end for;
end CFG_RAM512X18_VITAL;

---- CELL FIFO4K18 ----

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;
 
-- entity declaration --
entity FIFO4K18 is
  generic(
      TimingChecksOn   : Boolean := True;
      InstancePath     : String  := "*";
      Xon              : Boolean := False;
      MsgOn            : Boolean := True;
      
      tipd_AEVAL11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL10     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL9      : VitalDelayType01 := (0.000 ns, 0.000 ns);   	
      tipd_AEVAL8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL7      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL6      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL5      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL4      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL3      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL2      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AEVAL1      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AEVAL0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AFVAL11     : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AFVAL10     : VitalDelayType01 := (0.000 ns, 0.000 ns);      
      tipd_AFVAL9      : VitalDelayType01 := (0.000 ns, 0.000 ns);   
      tipd_AFVAL8      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_AFVAL7      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL6      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL5      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL4      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL3      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL2      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL1      : VitalDelayType01 := (0.000 ns, 0.000 ns); 
      tipd_AFVAL0      : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_REN         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RCLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RBLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WEN         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WBLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WCLK        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RESET       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RPIPE       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW2         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW1         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_RW0         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW2         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW1         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WW0         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_ESTOP       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_FSTOP       : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD17        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD16        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD15        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD14        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD13        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD12        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD11        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD10        : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD9         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD8         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD7         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD6         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD5         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD4         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD3         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD2         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD1         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_WD0         : VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_RCLK_RD17    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RCLK_RD16    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD15    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD14    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RCLK_RD13    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD12    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD11    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD10    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD9     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD8     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD7     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD6     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD5     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD4     : VitalDelayType01 := (0.100 ns, 0.100 ns);          
      tpd_RCLK_RD3     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD2     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD1     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_RD0     : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_EMPTY   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_AEMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RCLK_AFULL   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_WCLK_FULL    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_WCLK_AFULL   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_WCLK_AEMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD17   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD16   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD15   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD14   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD13   : VitalDelayType01 := (0.100 ns, 0.100 ns);          
      tpd_RESET_RD12   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD11   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD10   : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD9    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD8    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD7    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD6    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD5    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD4    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_RD3    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD2    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD1    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_RD0    : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_EMPTY  : VitalDelayType01 := (0.100 ns, 0.100 ns); 
      tpd_RESET_AEMPTY : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_FULL   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_RESET_AFULL  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tsetup_WD17_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD17_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD16_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD16_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD15_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD15_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD14_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD14_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD13_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD13_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD12_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD12_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD11_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD11_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD10_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD10_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WD9_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD9_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD8_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD8_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD7_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD7_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD6_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD6_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD5_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD5_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD4_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD4_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD3_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD3_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD2_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD2_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD1_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD1_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD0_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WD0_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD17_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD17_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD16_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD16_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD15_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD15_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD14_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD14_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD13_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD13_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD12_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD12_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD11_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD11_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD10_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD10_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WD9_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD9_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD8_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD8_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD7_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD7_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD6_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD6_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD5_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD5_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD4_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD4_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD3_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD3_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD2_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD2_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD1_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD1_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD0_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WD0_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      tsetup_WEN_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WEN_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WBLK_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WBLK_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_WEN_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WEN_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WBLK_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WBLK_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_REN_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_REN_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_RBLK_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_RBLK_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_REN_RCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_REN_RCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_RBLK_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      thold_RBLK_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_FSTOP_WCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_FSTOP_WCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_ESTOP_RCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      tsetup_ESTOP_RCLK_negedge_posedge    : VitalDelayType := 0.000 ns;
      thold_FSTOP_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_FSTOP_WCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      thold_ESTOP_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_ESTOP_RCLK_negedge_posedge     : VitalDelayType := 0.000 ns;
      tsetup_WW2_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WW2_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WW1_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WW1_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WW0_WCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_WW0_WCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_WW2_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WW2_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WW1_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WW1_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WW0_WCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_WW0_WCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      tsetup_RW2_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_RW2_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_RW1_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_RW1_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_RW0_RCLK_posedge_posedge      : VitalDelayType := 0.000 ns;
      tsetup_RW0_RCLK_negedge_posedge      : VitalDelayType := 0.000 ns;
      thold_RW2_RCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_RW2_RCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_RW1_RCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_RW1_RCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      thold_RW0_RCLK_posedge_posedge       : VitalDelayType := 0.000 ns;
      thold_RW0_RCLK_negedge_posedge       : VitalDelayType := 0.000 ns;
      tpw_WCLK_posedge                     : VitalDelayType := 0.000 ns;
      tpw_WCLK_negedge                     : VitalDelayType := 0.000 ns;
      tperiod_WCLK                         : VitalDelayType := 0.000 ns;                                     
      tpw_RCLK_posedge                     : VitalDelayType := 0.000 ns;                                   
      tpw_RCLK_negedge                     : VitalDelayType := 0.000 ns; 
      tperiod_RCLK                         : VitalDelayType := 0.000 ns;
      trecovery_RESET_RCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      trecovery_RESET_WCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_RESET_RCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      thold_RESET_WCLK_posedge_posedge     : VitalDelayType := 0.000 ns;
      tpw_RESET_negedge                    : VitalDelayType := 0.000 ns
     );

    port (
          AEVAL11	: IN STD_ULOGIC ;
          AEVAL10	: IN STD_ULOGIC ;
          AEVAL9	: IN STD_ULOGIC ;
          AEVAL8	: IN STD_ULOGIC ;
          AEVAL7	: IN STD_ULOGIC ;
          AEVAL6	: IN STD_ULOGIC ;
          AEVAL5	: IN STD_ULOGIC ;
          AEVAL4	: IN STD_ULOGIC ;
          AEVAL3	: IN STD_ULOGIC ;
          AEVAL2	: IN STD_ULOGIC ;
          AEVAL1	: IN STD_ULOGIC ;
          AEVAL0	: IN STD_ULOGIC ;
          AFVAL11	: IN STD_ULOGIC ;
          AFVAL10	: IN STD_ULOGIC ; 
          AFVAL9	: IN STD_ULOGIC ;
          AFVAL8	: IN STD_ULOGIC ;
          AFVAL7	: IN STD_ULOGIC ;
          AFVAL6	: IN STD_ULOGIC ;
          AFVAL5	: IN STD_ULOGIC ;
          AFVAL4	: IN STD_ULOGIC ;
          AFVAL3	: IN STD_ULOGIC ;
          AFVAL2	: IN STD_ULOGIC ;
          AFVAL1	: IN STD_ULOGIC ;
          AFVAL0	: IN STD_ULOGIC ;
          REN		: IN STD_ULOGIC ;
          RBLK		: IN STD_ULOGIC ;
          RCLK		: IN STD_ULOGIC ; 
          RESET		: IN STD_ULOGIC ;
          RPIPE		: IN STD_ULOGIC ;
          WEN		: IN STD_ULOGIC ;
          WBLK		: IN STD_ULOGIC ;
          WCLK		: IN STD_ULOGIC ;
          RW2		: IN STD_ULOGIC ;
          RW1		: IN STD_ULOGIC ;
          RW0		: IN STD_ULOGIC ;
          WW2		: IN STD_ULOGIC ;
          WW1		: IN STD_ULOGIC ;
          WW0		: IN STD_ULOGIC ;
          ESTOP		: IN STD_ULOGIC ;
          FSTOP		: IN STD_ULOGIC ;
          WD17		: IN STD_ULOGIC ;
          WD16		: IN STD_ULOGIC ;
          WD15		: IN STD_ULOGIC ;
          WD14		: IN STD_ULOGIC ;
          WD13		: IN STD_ULOGIC ;
          WD12		: IN STD_ULOGIC ;
          WD11		: IN STD_ULOGIC ;
          WD10		: IN STD_ULOGIC ;
          WD9		: IN STD_ULOGIC ;
          WD8		: IN STD_ULOGIC ;
          WD7		: IN STD_ULOGIC ;
          WD6		: IN STD_ULOGIC ;
          WD5		: IN STD_ULOGIC ;
          WD4		: IN STD_ULOGIC ;
          WD3		: IN STD_ULOGIC ;
          WD2		: IN STD_ULOGIC ;
          WD1		: IN STD_ULOGIC ;
          WD0		: IN STD_ULOGIC ;
          RD17		: OUT STD_ULOGIC ;
          RD16		: OUT STD_ULOGIC ;
          RD15		: OUT STD_ULOGIC ;
          RD14		: OUT STD_ULOGIC ;
          RD13		: OUT STD_ULOGIC ;
          RD12		: OUT STD_ULOGIC ;
          RD11		: OUT STD_ULOGIC ;
          RD10		: OUT STD_ULOGIC ;
          RD9		: OUT STD_ULOGIC ;
          RD8		: OUT STD_ULOGIC ;
          RD7		: OUT STD_ULOGIC ;
          RD6		: OUT STD_ULOGIC ; 
          RD5		: OUT STD_ULOGIC ;
          RD4		: OUT STD_ULOGIC ;
          RD3		: OUT STD_ULOGIC ;
          RD2		: OUT STD_ULOGIC ;
          RD1		: OUT STD_ULOGIC ;
          RD0		: OUT STD_ULOGIC ;
          FULL		: OUT STD_ULOGIC ;
          AFULL		: OUT STD_ULOGIC ;
          EMPTY		: OUT STD_ULOGIC ;
          AEMPTY	: OUT STD_ULOGIC 
         );  

   attribute VITAL_LEVEL0 of FIFO4K18 : entity is TRUE;

end FIFO4K18;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of FIFO4K18 is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal AFVAL11_ipd       : std_ulogic := 'X';
  signal AFVAL10_ipd       : std_ulogic := 'X';
  signal AFVAL9_ipd        : std_ulogic := 'X';
  signal AFVAL8_ipd        : std_ulogic := 'X';
  signal AFVAL7_ipd        : std_ulogic := 'X';
  signal AFVAL6_ipd        : std_ulogic := 'X';
  signal AFVAL5_ipd        : std_ulogic := 'X';
  signal AFVAL4_ipd        : std_ulogic := 'X';
  signal AFVAL3_ipd        : std_ulogic := 'X';
  signal AFVAL2_ipd        : std_ulogic := 'X';
  signal AFVAL1_ipd        : std_ulogic := 'X';
  signal AFVAL0_ipd        : std_ulogic := 'X';
  signal AEVAL11_ipd       : std_ulogic := 'X';
  signal AEVAL10_ipd       : std_ulogic := 'X'; 
  signal AEVAL9_ipd        : std_ulogic := 'X';
  signal AEVAL8_ipd        : std_ulogic := 'X';
  signal AEVAL7_ipd        : std_ulogic := 'X';
  signal AEVAL6_ipd        : std_ulogic := 'X';
  signal AEVAL5_ipd        : std_ulogic := 'X';
  signal AEVAL4_ipd        : std_ulogic := 'X';
  signal AEVAL3_ipd        : std_ulogic := 'X';
  signal AEVAL2_ipd        : std_ulogic := 'X';
  signal AEVAL1_ipd        : std_ulogic := 'X';
  signal AEVAL0_ipd        : std_ulogic := 'X';
  signal REN_ipd           : std_ulogic := 'X'; 
  signal RBLK_ipd          : std_ulogic := 'X'; 
  signal RCLK_ipd          : std_ulogic := 'X'; 
  signal RESET_ipd         : std_ulogic := 'X'; 
  signal RPIPE_ipd         : std_ulogic := 'X'; 
  signal WEN_ipd           : std_ulogic := 'X'; 
  signal WBLK_ipd          : std_ulogic := 'X'; 
  signal WCLK_ipd          : std_ulogic := 'X'; 
  signal RW2_ipd           : std_ulogic := 'X'; 
  signal RW1_ipd           : std_ulogic := 'X'; 
  signal RW0_ipd           : std_ulogic := 'X'; 
  signal WW2_ipd           : std_ulogic := 'X'; 
  signal WW1_ipd           : std_ulogic := 'X'; 
  signal WW0_ipd           : std_ulogic := 'X'; 
  signal ESTOP_ipd         : std_ulogic := 'X'; 
  signal FSTOP_ipd         : std_ulogic := 'X'; 
  signal WD17_ipd          : std_ulogic := 'X'; 
  signal WD16_ipd          : std_ulogic := 'X'; 
  signal WD15_ipd          : std_ulogic := 'X';  
  signal WD14_ipd          : std_ulogic := 'X'; 
  signal WD13_ipd          : std_ulogic := 'X'; 
  signal WD12_ipd          : std_ulogic := 'X'; 
  signal WD11_ipd          : std_ulogic := 'X'; 
  signal WD10_ipd          : std_ulogic := 'X'; 
  signal WD9_ipd           : std_ulogic := 'X'; 
  signal WD8_ipd           : std_ulogic := 'X'; 
  signal WD7_ipd           : std_ulogic := 'X'; 
  signal WD6_ipd           : std_ulogic := 'X'; 
  signal WD5_ipd           : std_ulogic := 'X'; 
  signal WD4_ipd           : std_ulogic := 'X'; 
  signal WD3_ipd           : std_ulogic := 'X'; 
  signal WD2_ipd           : std_ulogic := 'X'; 
  signal WD1_ipd           : std_ulogic := 'X'; 
  signal WD0_ipd           : std_ulogic := 'X';
  type MEM  is array(0 to 4095) of std_ulogic; -- Internal memory
  type MEM9 is array(0 to 511)  of std_ulogic; -- Internal memory


-- #########################################################
-- # Functions and Procedures
-- #########################################################

 FUNCTION get_max_address(width : integer) RETURN integer is
 variable max_address : integer := 0;
 BEGIN
     case width is
       when 1  =>  max_address := 4096;
       when 2  =>  max_address := 2048;
       when 4  =>  max_address := 1024;
       when 9  =>  max_address := 512;
       when 18 =>  max_address := 256;
       when others =>
                      assert false
                      report "Illegal width configuration"
                      severity Warning;
     end case;

     RETURN  max_address;
 end get_max_address;


 PROCEDURE increment_address_counter (
             variable ADDR        : INOUT integer;    -- Read/Write address
             variable wrap        : INOUT bit;        -- Wrap-around flag - toggles between 0 and 1
             variable width       : IN    integer;
             variable flag        : IN    std_ulogic; -- Empty/Full flag
             variable stop        : IN    std_ulogic  -- Estop/Fstop
            ) is

  variable depth :integer;

  BEGIN

  depth := get_max_address(width);
  if (flag = '0') then
    if (ADDR < depth - 1 ) then 
      ADDR := ADDR + 1;
    else
      ADDR := (ADDR + 1) mod depth;
      wrap := not wrap;
    end if;
  elsif ((flag = '1') and (stop = '0')) then
    if (ADDR < depth - 1 ) then
      ADDR := ADDR + 1;
    else
      ADDR := (ADDR + 1) mod depth;
      wrap := not wrap;
    end if;
  end if;
 END increment_address_counter;


 PROCEDURE fifo_flags (
                        variable  EMPTY          : INOUT std_ulogic;
                        variable  AEMPTY         : INOUT std_ulogic;
                        variable  FULL           : INOUT std_ulogic;
                        variable  AFULL          : INOUT std_ulogic;
                        variable  RADDR          : IN integer;
                        variable  RADDR_P2       : IN integer;
                        variable  RADDR_wrap     : IN bit;
                        variable  RADDR_wrap_P2  : IN bit;
                        variable  WADDR          : IN integer;
                        variable  WADDR_P2       : IN integer;
                        variable  WADDR_wrap     : IN bit;
                        variable  WADDR_wrap_P2  : IN bit;
                        variable  AFVAL          : IN integer;
                        variable  AEVAL          : IN integer;
                        variable  MAX_DEPTH      : IN integer;
                        variable  wwidth         : IN integer;
                        variable  rwidth         : IN integer;
                        variable  wwidth_bit     : IN integer;
                        variable  rwidth_bit     : IN integer
                      ) is

      variable raddr_rel : integer;
      variable waddr_rel : integer;
      variable raddr_rel_p2 : integer;
      variable waddr_rel_p2 : integer;
      variable rel_depth : integer;
      variable aeval_rel : integer;
      variable afval_rel : integer;
      variable num_fifo_entries : integer;
   BEGIN

     -- Pipelined addresses used for FULL and EMPTY calculations
     if (wwidth_bit < 0) then
       assert false
         report "Illegal Write port width configuration"
         severity warning;
     elsif (rwidth_bit < 0) then
       assert false
         report "Illegal Read port width configuration"
         severity warning;
     elsif (wwidth_bit >= rwidth_bit) then
       raddr_rel := RADDR /(2 ** (wwidth_bit - rwidth_bit));
       raddr_rel_p2 := RADDR_P2 /(2 ** (wwidth_bit - rwidth_bit));
       waddr_rel := WADDR;
       waddr_rel_p2 := WADDR_P2;
       rel_depth := 2 ** (12 - wwidth_bit);
       aeval_rel := AEVAL/(2 ** wwidth_bit);
       afval_rel := AFVAL/(2 ** wwidth_bit);
     else
       waddr_rel := WADDR /(2 ** (rwidth_bit - wwidth_bit));
       waddr_rel_p2 := WADDR_P2 /(2 ** (rwidth_bit - wwidth_bit));
       raddr_rel := RADDR;
       raddr_rel_p2 := RADDR_P2;
       rel_depth := 2 ** (12 - rwidth_bit);
       aeval_rel := AEVAL/(2 ** rwidth_bit);
       afval_rel := AFVAL/(2 ** rwidth_bit);       
     end if;
    
     if ((WADDR_wrap = RADDR_wrap_P2) and ( waddr_rel = raddr_rel_p2 )) then
       FULL := '1';
     else
       FULL := '0';
     end if;

     if ((RADDR_wrap = WADDR_wrap_P2) and (waddr_rel_p2 = raddr_rel)) then
       EMPTY := '1';
     else
       EMPTY := '0';
     end if;
     
     -- Number of FIFO ENTRIES
     if (waddr_rel >= raddr_rel) then
       num_fifo_entries := waddr_rel - raddr_rel;
     else
       num_fifo_entries := rel_depth + waddr_rel - raddr_rel;
     end if;
     --aempty, afull generation
     if (FULL = '1') then
       AEMPTY := '0';
     else
       if(aeval_rel >= 0) then
         if (num_fifo_entries > aeval_rel) then 
           AEMPTY := '0';
         else
           AEMPTY := '1';
         end if;
       end if;
     end if;

     if (EMPTY = '1') then
       AFULL := '0';
     elsif (FULL = '1') then
       AFULL := '1';
     else
       if(afval_rel >= 0) then 
         if (num_fifo_entries < afval_rel) then
           AFULL := '0';
         else
           AFULL := '1';
         end if;
       end if;
     end if;
     
 END fifo_flags;

 begin   --  VITAL_ACT

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WireDelay: block

  begin --  block WireDelay
    VitalWireDelay (AEVAL11_ipd, AEVAL11, VitalExtendToFillDelay(tipd_AEVAL11));
    VitalWireDelay (AEVAL10_ipd, AEVAL10, VitalExtendToFillDelay(tipd_AEVAL10));
    VitalWireDelay (AEVAL9_ipd, AEVAL9, VitalExtendToFillDelay(tipd_AEVAL9));
    VitalWireDelay (AEVAL8_ipd, AEVAL8, VitalExtendToFillDelay(tipd_AEVAL8));
    VitalWireDelay (AEVAL7_ipd, AEVAL7, VitalExtendToFillDelay(tipd_AEVAL7));
    VitalWireDelay (AEVAL6_ipd, AEVAL6, VitalExtendToFillDelay(tipd_AEVAL6));
    VitalWireDelay (AEVAL5_ipd, AEVAL5, VitalExtendToFillDelay(tipd_AEVAL5));
    VitalWireDelay (AEVAL4_ipd, AEVAL4, VitalExtendToFillDelay(tipd_AEVAL4));
    VitalWireDelay (AEVAL3_ipd, AEVAL3, VitalExtendToFillDelay(tipd_AEVAL3));
    VitalWireDelay (AEVAL2_ipd, AEVAL2, VitalExtendToFillDelay(tipd_AEVAL2));
    VitalWireDelay (AEVAL1_ipd, AEVAL1, VitalExtendToFillDelay(tipd_AEVAL1));
    VitalWireDelay (AEVAL0_ipd, AEVAL0, VitalExtendToFillDelay(tipd_AEVAL0));
    VitalWireDelay (AFVAL11_ipd, AFVAL11, VitalExtendToFillDelay(tipd_AFVAL11));
    VitalWireDelay (AFVAL10_ipd, AFVAL10, VitalExtendToFillDelay(tipd_AFVAL10));
    VitalWireDelay (AFVAL9_ipd, AFVAL9, VitalExtendToFillDelay(tipd_AFVAL9));
    VitalWireDelay (AFVAL8_ipd, AFVAL8, VitalExtendToFillDelay(tipd_AFVAL8));
    VitalWireDelay (AFVAL7_ipd, AFVAL7, VitalExtendToFillDelay(tipd_AFVAL7));
    VitalWireDelay (AFVAL6_ipd, AFVAL6, VitalExtendToFillDelay(tipd_AFVAL6));
    VitalWireDelay (AFVAL5_ipd, AFVAL5, VitalExtendToFillDelay(tipd_AFVAL5));
    VitalWireDelay (AFVAL4_ipd, AFVAL4, VitalExtendToFillDelay(tipd_AFVAL4));
    VitalWireDelay (AFVAL3_ipd, AFVAL3, VitalExtendToFillDelay(tipd_AFVAL3));
    VitalWireDelay (AFVAL2_ipd, AFVAL2, VitalExtendToFillDelay(tipd_AFVAL2));
    VitalWireDelay (AFVAL1_ipd, AFVAL1, VitalExtendToFillDelay(tipd_AFVAL1));
    VitalWireDelay (AFVAL0_ipd, AFVAL0, VitalExtendToFillDelay(tipd_AFVAL0));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN)); 
    VitalWireDelay (RBLK_ipd, RBLK, VitalExtendToFillDelay(tipd_RBLK));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK)); 
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN)); 
    VitalWireDelay (WBLK_ipd, WBLK, VitalExtendToFillDelay(tipd_WBLK));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET)); 
    VitalWireDelay (RPIPE_ipd, RPIPE, VitalExtendToFillDelay(tipd_RPIPE));
    VitalWireDelay (RW2_ipd, RW2, VitalExtendToFillDelay(tipd_RW2)); 
    VitalWireDelay (RW1_ipd, RW1, VitalExtendToFillDelay(tipd_RW1)); 
    VitalWireDelay (RW0_ipd, RW0, VitalExtendToFillDelay(tipd_RW0)); 
    VitalWireDelay (WW2_ipd, WW2, VitalExtendToFillDelay(tipd_WW2)); 
    VitalWireDelay (WW1_ipd, WW1, VitalExtendToFillDelay(tipd_WW1)); 
    VitalWireDelay (WW0_ipd, WW0, VitalExtendToFillDelay(tipd_WW0)); 
    VitalWireDelay (ESTOP_ipd, ESTOP, VitalExtendToFillDelay(tipd_ESTOP)); 
    VitalWireDelay (FSTOP_ipd, FSTOP, VitalExtendToFillDelay(tipd_FSTOP)); 
    VitalWireDelay (WD17_ipd, WD17, VitalExtendToFillDelay(tipd_WD17));  
    VitalWireDelay (WD16_ipd, WD16, VitalExtendToFillDelay(tipd_WD16));
    VitalWireDelay (WD15_ipd, WD15, VitalExtendToFillDelay(tipd_WD15));
    VitalWireDelay (WD14_ipd, WD14, VitalExtendToFillDelay(tipd_WD14));
    VitalWireDelay (WD13_ipd, WD13, VitalExtendToFillDelay(tipd_WD13));
    VitalWireDelay (WD12_ipd, WD12, VitalExtendToFillDelay(tipd_WD12));
    VitalWireDelay (WD11_ipd, WD11, VitalExtendToFillDelay(tipd_WD11));
    VitalWireDelay (WD10_ipd, WD10, VitalExtendToFillDelay(tipd_WD10));
    VitalWireDelay (WD9_ipd, WD9, VitalExtendToFillDelay(tipd_WD9));
    VitalWireDelay (WD8_ipd, WD8, VitalExtendToFillDelay(tipd_WD8));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0)); 


   end block WireDelay;


  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (AEVAL11_ipd, AEVAL10_ipd, AEVAL9_ipd, AEVAL8_ipd, AEVAL7_ipd, 
                           AEVAL6_ipd, AEVAL5_ipd, AEVAL4_ipd, AEVAL3_ipd, AEVAL2_ipd,
                           AEVAL1_ipd, AEVAL0_ipd, AFVAL11_ipd, AFVAL10_ipd, AFVAL9_ipd,
                           AFVAL8_ipd, AFVAL7_ipd, AFVAL6_ipd, AFVAL5_ipd, AFVAL4_ipd,
                           AFVAL3_ipd, AFVAL2_ipd, AFVAL1_ipd, AFVAL0_ipd, REN_ipd, 
                           RBLK_ipd, RCLK_ipd, WEN_ipd, WBLK_ipd, WCLK_ipd, RESET_ipd,
                           RPIPE_ipd, RW2_ipd, RW1_ipd, RW0_ipd, WW2_ipd, WW1_ipd,
                           WW0_ipd, ESTOP_ipd, FSTOP_ipd, WD17_ipd, WD16_ipd, WD15_ipd,
                           WD14_ipd, WD13_ipd, WD12_ipd, WD11_ipd, WD10_ipd, WD9_ipd,
                           WD8_ipd, WD7_ipd, WD6_ipd, WD5_ipd, WD4_ipd, WD3_ipd, WD2_ipd,
                           WD1_ipd, WD0_ipd)

  -- some internal veriable declaration
     variable afullvalue    : integer := 0;
     variable aemptyvalue   : integer := 0;
     variable WADDR         : integer;-- := 0;
     variable WADDR_P1      : integer;-- := 0;
     variable WADDR_P2      : integer;-- := 0;
     variable WADDR_wrap    : bit   ;--  := '0';
     variable WADDR_wrap_P1 : bit   ;--  := '0';
     variable WADDR_wrap_P2 : bit   ;--  := '0';
     variable RADDR         : integer;-- := 0;
     variable RADDR_P1      : integer;-- := 0;
     variable RADDR_P2      : integer;-- := 0;
     variable RADDR_wrap    : bit    ;-- := '0';
     variable RADDR_wrap_P1 : bit    ;-- := '1';
     variable RADDR_wrap_P2 : bit    ;-- := '1';

     variable wwidth        : integer;
     variable rwidth        : integer;
     variable wwidth_bit        : integer;
     variable rwidth_bit        : integer;
     variable rmask : std_ulogic_vector(3 downto 0);
     variable wmask : std_ulogic_vector(3 downto 0);
     variable mask : std_ulogic_vector(3 downto 0);
     variable MAX_depth     : integer := 4095;
     variable MEM_TMP       : MEM;
     variable MEM9_TMP      : MEM9;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-4095, -4095, 0, 1, -4095, -4095, 0, 1, -4095);

     
     --  Read Timing Check Results
     variable Tviol_WD17_WCLK_posedge : X01 := '0';
     variable TmDt_WD17_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD16_WCLK_posedge : X01 := '0';
     variable TmDt_WD16_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD15_WCLK_posedge : X01 := '0';
     variable TmDt_WD15_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD14_WCLK_posedge : X01 := '0';
     variable TmDt_WD14_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD13_WCLK_posedge : X01 := '0';
     variable TmDt_WD13_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD12_WCLK_posedge : X01 := '0';
     variable TmDt_WD12_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD11_WCLK_posedge : X01 := '0';
     variable TmDt_WD11_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD10_WCLK_posedge : X01 := '0';
     variable TmDt_WD10_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD9_WCLK_posedge : X01 := '0';
     variable TmDt_WD9_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD8_WCLK_posedge : X01 := '0';
     variable TmDt_WD8_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLK_WCLK_posedge : X01 := '0';
     variable TmDt_WBLK_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_FSTOP_WCLK_posedge : X01 := '0';
     variable TmDt_FSTOP_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLK_RCLK_posedge : X01 := '0';
     variable TmDt_RBLK_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_ESTOP_RCLK_posedge : X01 := '0';
     variable TmDt_ESTOP_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW2_WCLK_posedge : X01 := '0';
     variable TmDt_WW2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW1_WCLK_posedge : X01 := '0';
     variable TmDt_WW1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WW0_WCLK_posedge : X01 := '0';
     variable TmDt_WW0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW2_RCLK_posedge : X01 := '0';
     variable TmDt_RW2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW1_RCLK_posedge : X01 := '0';
     variable TmDt_RW1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RW0_RCLK_posedge : X01 := '0';
     variable TmDt_RW0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;

     
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
     variable Tviol_RESET_RCLK_posedge : X01 := '0';
     variable Tmkr_RESET_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLK_posedge : X01 := '0';
     variable Tmkr_RESET_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RESET : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET : X01 := '0';

    
   -- functional Results

     variable RD0_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD7_zd : std_ulogic;
     variable RD8_zd : std_ulogic;
     variable RD9_zd : std_ulogic;
     variable RD10_zd : std_ulogic;
     variable RD11_zd : std_ulogic;
     variable RD12_zd : std_ulogic;
     variable RD13_zd : std_ulogic;
     variable RD14_zd : std_ulogic;
     variable RD15_zd : std_ulogic;
     variable RD16_zd : std_ulogic;
     variable RD17_zd : std_ulogic;
     variable FULL_zd : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable AFULL_zd : std_ulogic;
     variable AEMPTY_zd : std_ulogic; 

     variable RD0_stg : std_ulogic;
     variable RD1_stg : std_ulogic;
     variable RD2_stg : std_ulogic;
     variable RD3_stg : std_ulogic;
     variable RD4_stg : std_ulogic;
     variable RD5_stg : std_ulogic;
     variable RD6_stg : std_ulogic;
     variable RD7_stg : std_ulogic;
     variable RD8_stg : std_ulogic;
     variable RD9_stg : std_ulogic;
     variable RD10_stg : std_ulogic;
     variable RD11_stg : std_ulogic;
     variable RD12_stg : std_ulogic;
     variable RD13_stg : std_ulogic;
     variable RD14_stg : std_ulogic;
     variable RD15_stg : std_ulogic;
     variable RD16_stg : std_ulogic;
     variable RD17_stg : std_ulogic;

   -- Output Glitch Detection Support Variables

     variable RD0_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD8_GlitchData : VitalGlitchDataType;
     variable RD9_GlitchData : VitalGlitchDataType;
     variable RD10_GlitchData : VitalGlitchDataType;
     variable RD11_GlitchData : VitalGlitchDataType;
     variable RD12_GlitchData : VitalGlitchDataType;
     variable RD13_GlitchData : VitalGlitchDataType;
     variable RD14_GlitchData : VitalGlitchDataType;
     variable RD15_GlitchData : VitalGlitchDataType;
     variable RD16_GlitchData : VitalGlitchDataType;
     variable RD17_GlitchData : VitalGlitchDataType;
     variable FULL_GlitchData : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable AFULL_GlitchData : VitalGlitchDataType;
     variable AEMPTY_GlitchData : VitalGlitchDataType;
    
       -- last value variables
     variable WCLK_previous : std_ulogic := '0';
     variable RCLK_previous : std_ulogic := '0';
 
     variable issue_WBLK : std_ulogic := '0';
     variable issue_WEN : std_ulogic := '0';
     variable issue_RBLK : std_ulogic := '0';
     variable issue_REN : std_ulogic := '0';
     variable issue_FSTOP : std_ulogic := '0';
     variable issue_ESTOP : std_ulogic := '0';
     variable issue_AFVAL : std_ulogic := '0';     
     variable issue_AEVAL : std_ulogic := '0';     

     variable RPIPE_delayed : std_ulogic := 'X';
     variable RESET_delayed : std_ulogic := 'X';
     variable WD0_delayed  : std_ulogic := 'X';
     variable WD1_delayed  : std_ulogic := 'X';
     variable WD2_delayed  : std_ulogic := 'X';
     variable WD3_delayed  : std_ulogic := 'X';
     variable WD4_delayed  : std_ulogic := 'X';
     variable WD5_delayed  : std_ulogic := 'X';
     variable WD6_delayed  : std_ulogic := 'X';
     variable WD7_delayed  : std_ulogic := 'X';
     variable WD8_delayed  : std_ulogic := 'X';
     variable WD9_delayed  : std_ulogic := 'X';
     variable WD10_delayed  : std_ulogic := 'X';
     variable WD11_delayed  : std_ulogic := 'X';
     variable WD12_delayed  : std_ulogic := 'X';
     variable WD13_delayed  : std_ulogic := 'X';
     variable WD14_delayed  : std_ulogic := 'X';
     variable WD15_delayed  : std_ulogic := 'X';
     variable WD16_delayed  : std_ulogic := 'X';
     variable WD17_delayed  : std_ulogic := 'X';
     variable ESTOP_delayed : std_ulogic := 'X';
     variable FSTOP_delayed : std_ulogic := 'X';
 
 begin -- process VITALBehavior

if (TimingChecksOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------
   
 -- setup / hold check for RCLK to RESET signal ;
       VitalSetupHoldCheck ( Tviol_RESET_RCLK_posedge,
                             Tmkr_RESET_RCLK_posedge,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             trecovery_RESET_RCLK_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_RESET_RCLK_posedge_posedge,
                             (TO_X01(REN_ipd) = '1') and (TO_X01(RBLK_ipd) = '0'),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

  -- setup / hold check for WCLK to RESET signal ;
       VitalSetupHoldCheck ( Tviol_RESET_WCLK_posedge,
                             Tmkr_RESET_WCLK_posedge,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             trecovery_RESET_WCLK_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_RESET_WCLK_posedge_posedge,
                             (TO_X01(WEN_ipd) = '1') and (TO_X01(WBLK_ipd) = '0'),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                             TmDt_REN_RCLK_posedge,
                             REN_ipd, "REN",
                             0.0 ns,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                         tsetup_REN_RCLK_posedge_posedge,
                         tsetup_REN_RCLK_negedge_posedge,
                         thold_REN_RCLK_posedge_posedge,
                         thold_REN_RCLK_negedge_posedge,
                             ((TO_X01(RBLK_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLK_RCLK_posedge,
                             TmDt_RBLK_RCLK_posedge,
                             RBLK_ipd, "RBLK",
                             0.0 ns,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                         tsetup_RBLK_RCLK_posedge_posedge,
                         tsetup_RBLK_RCLK_negedge_posedge,
                         thold_RBLK_RCLK_posedge_posedge,
                         thold_RBLK_RCLK_negedge_posedge,
                             ((TO_X01(REN_ipd) = '1') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

      -- setup hold WEN, WBLK low when WCLK rising
       VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                             TmDt_WEN_WCLK_posedge,
                             WEN_ipd, "WEN",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_WEN_WCLK_posedge_posedge,
                         tsetup_WEN_WCLK_negedge_posedge,
                         thold_WEN_WCLK_posedge_posedge,
                         thold_WEN_WCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLK_WCLK_posedge,
                             TmDt_WBLK_WCLK_posedge,
                             WBLK_ipd, "WBLK",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_WBLK_WCLK_posedge_posedge,
                         tsetup_WBLK_WCLK_negedge_posedge,
                         thold_WBLK_WCLK_posedge_posedge,
                         thold_WBLK_WCLK_negedge_posedge,
                             ((TO_X01(WEN_ipd) = '1') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       -- setup hold FSTOP when WCLK rising
       VitalSetupHoldCheck ( Tviol_FSTOP_WCLK_posedge,
                             TmDt_FSTOP_WCLK_posedge,
                             FSTOP_ipd, "FSTOP",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_FSTOP_WCLK_posedge_posedge,
                         tsetup_FSTOP_WCLK_negedge_posedge,
                         thold_FSTOP_WCLK_posedge_posedge,
                         thold_FSTOP_WCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );
         -- setup hold ESTOP when RCLK rising
       VitalSetupHoldCheck ( Tviol_ESTOP_RCLK_posedge,
                             TmDt_ESTOP_RCLK_posedge,
                             ESTOP_ipd, "ESTOP",
                             0.0 ns,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                         tsetup_ESTOP_RCLK_posedge_posedge,
                         tsetup_ESTOP_RCLK_negedge_posedge,
                         thold_ESTOP_RCLK_posedge_posedge,
                         thold_ESTOP_RCLK_negedge_posedge,
                             ((TO_X01(RBLK_ipd) = '0') and (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );


         -- setup hold WW2,WW1,WW0 when WCLK rising
       VitalSetupHoldCheck ( Tviol_WW2_WCLK_posedge,
                             TmDt_WW2_WCLK_posedge,
                             WW2_ipd, "WW2",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_WW2_WCLK_posedge_posedge,
                         tsetup_WW2_WCLK_negedge_posedge,
                         thold_WW2_WCLK_posedge_posedge,
                         thold_WW2_WCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WW1_WCLK_posedge,
                             TmDt_WW1_WCLK_posedge,
                             WW1_ipd, "WW1",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_WW1_WCLK_posedge_posedge,
                         tsetup_WW1_WCLK_negedge_posedge,
                         thold_WW1_WCLK_posedge_posedge,
                         thold_WW1_WCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WW0_WCLK_posedge,
                             TmDt_WW0_WCLK_posedge,
                             WW0_ipd, "WW0",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_WW0_WCLK_posedge_posedge,
                         tsetup_WW0_WCLK_negedge_posedge,
                         thold_WW0_WCLK_posedge_posedge,
                         thold_WW0_WCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

      
        -- setup hold RW2,RW1,RW0 when RCLK rising
       VitalSetupHoldCheck ( Tviol_RW2_RCLK_posedge,
                             TmDt_RW2_RCLK_posedge,
                             RW2_ipd, "RW2",
                             0.0 ns,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                         tsetup_RW2_RCLK_posedge_posedge,
                         tsetup_RW2_RCLK_negedge_posedge,
                         thold_RW2_RCLK_posedge_posedge,
                         thold_RW2_RCLK_negedge_posedge,
                             ((TO_X01(RBLK_ipd) = '0') and (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RW1_RCLK_posedge,
                             TmDt_RW1_RCLK_posedge,
                             RW1_ipd, "RW1",
                             0.0 ns,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                         tsetup_RW1_RCLK_posedge_posedge,
                         tsetup_RW1_RCLK_negedge_posedge,
                         thold_RW1_RCLK_posedge_posedge,
                         thold_RW1_RCLK_negedge_posedge,
                             ((TO_X01(RBLK_ipd) = '0') and (TO_X01(REN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_RW0_RCLK_posedge,
                             TmDt_RW0_RCLK_posedge,
                             RW0_ipd, "RW0",
                             0.0 ns,
                             RCLK_ipd, "RCLK",
                             0.0 ns,
                         tsetup_RW0_RCLK_posedge_posedge,
                         tsetup_RW0_RCLK_negedge_posedge,
                         thold_RW0_RCLK_posedge_posedge,
                         thold_RW0_RCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

              -- setup hold WD17-0 when WCLK rising
              VitalSetupHoldCheck ( Tviol_WD17_WCLK_posedge,
                             TmDt_WD17_WCLK_posedge,
                             WD17_ipd, "WD17",
                             0.0 ns,
                             WCLK_ipd, "WCLK",
                             0.0 ns,
                         tsetup_WD17_WCLK_posedge_posedge,
                         tsetup_WD17_WCLK_negedge_posedge,
                         thold_WD17_WCLK_posedge_posedge,
                         thold_WD17_WCLK_negedge_posedge,
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/ FIFO4K18",
                             TRUE,
                             TRUE,
                             WARNING
                             );

               VitalSetupHoldCheck ( Tviol_WD16_WCLK_posedge,           
                             TmDt_WD16_WCLK_posedge,            
                             WD16_ipd, "WD16",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD16_WCLK_posedge_posedge,          
                         tsetup_WD16_WCLK_negedge_posedge,          
                         thold_WD16_WCLK_posedge_posedge,           
                         thold_WD16_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
               VitalSetupHoldCheck ( Tviol_WD15_WCLK_posedge,           
                             TmDt_WD15_WCLK_posedge,            
                             WD15_ipd, "WD15",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD15_WCLK_posedge_posedge,          
                         tsetup_WD15_WCLK_negedge_posedge,          
                         thold_WD15_WCLK_posedge_posedge,           
                         thold_WD15_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
              VitalSetupHoldCheck ( Tviol_WD14_WCLK_posedge,           
                             TmDt_WD14_WCLK_posedge,            
                             WD14_ipd, "WD14",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD14_WCLK_posedge_posedge,          
                         tsetup_WD14_WCLK_negedge_posedge,          
                         thold_WD14_WCLK_posedge_posedge,           
                         thold_WD14_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
             VitalSetupHoldCheck ( Tviol_WD13_WCLK_posedge,           
                             TmDt_WD13_WCLK_posedge,            
                             WD13_ipd, "WD13",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD13_WCLK_posedge_posedge,          
                         tsetup_WD13_WCLK_negedge_posedge,          
                         thold_WD13_WCLK_posedge_posedge,           
                         thold_WD13_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
            VitalSetupHoldCheck ( Tviol_WD12_WCLK_posedge,           
                             TmDt_WD12_WCLK_posedge,            
                             WD12_ipd, "WD12",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD12_WCLK_posedge_posedge,          
                         tsetup_WD12_WCLK_negedge_posedge,          
                         thold_WD12_WCLK_posedge_posedge,           
                         thold_WD12_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
            VitalSetupHoldCheck ( Tviol_WD11_WCLK_posedge,           
                             TmDt_WD11_WCLK_posedge,            
                             WD11_ipd, "WD11",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD11_WCLK_posedge_posedge,          
                         tsetup_WD11_WCLK_negedge_posedge,          
                         thold_WD11_WCLK_posedge_posedge,           
                         thold_WD11_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
            VitalSetupHoldCheck ( Tviol_WD10_WCLK_posedge,           
                             TmDt_WD10_WCLK_posedge,            
                             WD10_ipd, "WD10",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD10_WCLK_posedge_posedge,          
                         tsetup_WD10_WCLK_negedge_posedge,          
                         thold_WD10_WCLK_posedge_posedge,           
                         thold_WD10_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
            VitalSetupHoldCheck ( Tviol_WD9_WCLK_posedge,           
                             TmDt_WD9_WCLK_posedge,            
                             WD9_ipd, "WD9",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD9_WCLK_posedge_posedge,          
                         tsetup_WD9_WCLK_negedge_posedge,          
                         thold_WD9_WCLK_posedge_posedge,           
                         thold_WD9_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
            VitalSetupHoldCheck ( Tviol_WD8_WCLK_posedge,           
                             TmDt_WD8_WCLK_posedge,            
                             WD8_ipd, "WD8",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD8_WCLK_posedge_posedge,          
                         tsetup_WD8_WCLK_negedge_posedge,          
                         thold_WD8_WCLK_posedge_posedge,           
                         thold_WD8_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
            VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,           
                             TmDt_WD7_WCLK_posedge,            
                             WD7_ipd, "WD7",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD7_WCLK_posedge_posedge,          
                         tsetup_WD7_WCLK_negedge_posedge,          
                         thold_WD7_WCLK_posedge_posedge,           
                         thold_WD7_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
           VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,           
                             TmDt_WD6_WCLK_posedge,            
                             WD6_ipd, "WD6",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD6_WCLK_posedge_posedge,          
                         tsetup_WD6_WCLK_negedge_posedge,          
                         thold_WD6_WCLK_posedge_posedge,           
                         thold_WD6_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
          VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,           
                             TmDt_WD5_WCLK_posedge,            
                             WD5_ipd, "WD5",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD5_WCLK_posedge_posedge,          
                         tsetup_WD5_WCLK_negedge_posedge,          
                         thold_WD5_WCLK_posedge_posedge,           
                         thold_WD5_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
         VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,           
                             TmDt_WD4_WCLK_posedge,            
                             WD4_ipd, "WD4",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD4_WCLK_posedge_posedge,          
                         tsetup_WD4_WCLK_negedge_posedge,          
                         thold_WD4_WCLK_posedge_posedge,           
                         thold_WD4_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
         VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,           
                             TmDt_WD3_WCLK_posedge,            
                             WD3_ipd, "WD3",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD3_WCLK_posedge_posedge,          
                         tsetup_WD3_WCLK_negedge_posedge,          
                         thold_WD3_WCLK_posedge_posedge,           
                         thold_WD3_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
         VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,           
                             TmDt_WD2_WCLK_posedge,            
                             WD2_ipd, "WD2",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD2_WCLK_posedge_posedge,          
                         tsetup_WD2_WCLK_negedge_posedge,          
                         thold_WD2_WCLK_posedge_posedge,           
                         thold_WD2_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
       VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,           
                             TmDt_WD1_WCLK_posedge,            
                             WD1_ipd, "WD1",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD1_WCLK_posedge_posedge,          
                         tsetup_WD1_WCLK_negedge_posedge,          
                         thold_WD1_WCLK_posedge_posedge,           
                         thold_WD1_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        
       VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,           
                             TmDt_WD0_WCLK_posedge,            
                             WD0_ipd, "WD0",           
                             0.0 ns,           
                             WCLK_ipd, "WCLK",         
                             0.0 ns,           
                         tsetup_WD0_WCLK_posedge_posedge,          
                         tsetup_WD0_WCLK_negedge_posedge,          
                         thold_WD0_WCLK_posedge_posedge,           
                         thold_WD0_WCLK_negedge_posedge,           
                             ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0') and (TO_X01(RESET_ipd) = '1')),             
                             '/',              
                             InstancePath & "/ FIFO4K18",              
                             TRUE,             
                             TRUE,             
                             WARNING           
                             );        


 --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLK,
                              PeriodData_RCLK,
                              RCLK_ipd, "RCLK",
                              0.0 ns,
                              tperiod_RCLK,
                              tpw_RCLK_posedge,
                              tpw_RCLK_negedge,
                              (TO_X01(REN_ipd) = '1') and (TO_X01(RBLK_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
                              InstancePath & "/ FIFO4K18",
                              TRUE,
                              TRUE,
                              WARNING
                              );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLK,
                              PeriodData_WCLK,
                              WCLK_ipd, "WCLK",
                              0.0 ns,
                              tperiod_WCLK,
                              tpw_WCLK_posedge,
                              tpw_WCLK_negedge,
                              (TO_X01(REN_ipd) = '1') and (TO_X01(RBLK_ipd) = '0') and (TO_X01(RESET_ipd) = '1'),
                              InstancePath & "/ FIFO4K18",
                              TRUE,
                              TRUE,
                              WARNING
                              );

  

      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              TRUE,
                              InstancePath & "/ FIFO4K18",
                              TRUE,
                              TRUE,
                              WARNING
                              );
     end if;

 
  if ((TO_X01(WW2_ipd) = '0') and (TO_X01(WW1_ipd) = '0') and (TO_X01(WW0_ipd) = '0')) then
    wwidth := 1;
    wwidth_bit := 0;
    wmask := "1111";
  elsif ((TO_X01(WW2_ipd) = '0') and (TO_X01(WW1_ipd) = '0') and (TO_X01(WW0_ipd) = '1')) then
    wwidth := 2;
    wwidth_bit := 1 ;
    wmask := "1110";
  elsif ((TO_X01(WW2_ipd) = '0') and (TO_X01(WW1_ipd) = '1') and (TO_X01(WW0_ipd) = '0')) then
    wwidth := 4;
     wwidth_bit := 2;
    wmask := "1100";
  elsif ((TO_X01(WW2_ipd) = '0') and (TO_X01(WW1_ipd) = '1') and (TO_X01(WW0_ipd) = '1')) then
    wwidth := 9;
     wwidth_bit := 3;
    wmask := "1000";
  elsif ((TO_X01(WW2_ipd) = '1') and (TO_X01(WW1_ipd) = '0') and (TO_X01(WW0_ipd) = '0')) then
    wwidth := 18;
     wwidth_bit := 4;
    wmask := "0000";
  else
    wwidth := -1;
     wwidth_bit := -1;
    wmask := "XXXX";
  end if;

  if ((TO_X01(RW2_ipd) = '0') and (TO_X01(RW1_ipd) = '0') and (TO_X01(RW0_ipd) = '0')) then
    rwidth := 1;
    rwidth_bit := 0;
    rmask := "1111";
  elsif ((TO_X01(RW2_ipd) = '0') and (TO_X01(RW1_ipd) = '0') and (TO_X01(RW0_ipd) = '1')) then
    rwidth := 2;
    rwidth_bit := 1;
    rmask := "1110";
  elsif ((TO_X01(RW2_ipd) = '0') and (TO_X01(RW1_ipd) = '1') and (TO_X01(RW0_ipd) = '0')) then
    rwidth := 4;
    rwidth_bit := 2;
    rmask := "1100";
  elsif ((TO_X01(RW2_ipd) = '0') and (TO_X01(RW1_ipd) = '1') and (TO_X01(RW0_ipd) = '1')) then
    rwidth := 9;
    rwidth_bit := 3;
    rmask := "1000";
  elsif ((TO_X01(RW2_ipd) = '1') and (TO_X01(RW1_ipd) = '0') and (TO_X01(RW0_ipd) = '0')) then
    rwidth := 18;
    rwidth_bit := 4;
    rmask := "0000";
  else
    rwidth := -1;
    rwidth_bit := -1;
    rmask := "XXXX";
  end if;

mask := rmask and wmask;

  -----------------------------------------------------------
  --    calculate the almost FULL and almost EMPTY value   --
  -----------------------------------------------------------

  afullvalue := ((INT(AFVAL11_ipd)*2048) + (INT(AFVAL10_ipd)*1024) +
                (INT(AFVAL9_ipd)*512)   + (INT(AFVAL8_ipd)*256)   +
                (INT(AFVAL7_ipd)*128)   + (INT(AFVAL6_ipd)*64)    +
                (INT(AFVAL5_ipd)*32)    + (INT(AFVAL4_ipd)*16)    +
                (INT(AFVAL3_ipd and mask(3))*8) +
                (INT(AFVAL2_ipd and mask(2))*4) +
                (INT(AFVAL1_ipd and mask(1))*2) +
                (INT(AFVAL0_ipd and mask(0))*1));

  aemptyvalue := ((INT(AEVAL11_ipd)*2048) + (INT(AEVAL10_ipd)*1024) +
                (INT(AEVAL9_ipd)*512)   + (INT(AEVAL8_ipd)*256)   +
                (INT(AEVAL7_ipd)*128)   + (INT(AEVAL6_ipd)*64)    +
                (INT(AEVAL5_ipd)*32)    + (INT(AEVAL4_ipd)*16)    +
                (INT(AEVAL3_ipd and mask(3))*8) +
                (INT(AEVAL2_ipd and mask(2))*4)     +
                (INT(AEVAL1_ipd and mask(1))*2)     +
                (INT(AEVAL0_ipd and mask(0))*1));



  ------------------------------------------------------------
  --               FIFO RESET                               --
  ------------------------------------------------------------
  
  if (TO_X01(RESET_ipd) = 'X') then
    if(RESET_ipd'event and TO_X01(RESET_ipd'last_value) /= 'X') then
      assert false
        report "RESET signal unknown."
        severity Warning;
    end if;
  elsif (TO_X01(RESET_ipd) = '0') then
    WADDR := 0;
    WADDR_P1 := 0;
    WADDR_P2 := 0;
    WADDR_wrap := '0';
    WADDR_wrap_P1 := '0';
    WADDR_wrap_P2 := '0';
    RADDR := 0;
    RADDR_P1 := 0;
    RADDR_P2 := 0;
    RADDR_wrap := '0';
    RADDR_wrap_P1 := '1';
    RADDR_wrap_P2 := '1';
    FULL_zd := '0';
    EMPTY_zd := '1';
    AFULL_zd := '0';
    AEMPTY_zd := '1';
    RD0_zd  := '0';
    RD1_zd  := '0';
    RD2_zd  := '0';
    RD3_zd  := '0';
    RD4_zd  := '0';
    RD5_zd  := '0';
    RD6_zd  := '0';
    RD7_zd  := '0';
    RD8_zd  := '0';
    RD9_zd  := '0'; 
    RD10_zd := '0'; 
    RD11_zd := '0'; 
    RD12_zd := '0'; 
    RD13_zd := '0'; 
    RD14_zd := '0'; 
    RD15_zd := '0'; 
    RD16_zd := '0'; 
    RD17_zd := '0';

    RD0_stg  := '0';
    RD1_stg  := '0';
    RD2_stg  := '0';
    RD3_stg  := '0';
    RD4_stg  := '0';
    RD5_stg  := '0';
    RD6_stg  := '0';
    RD7_stg  := '0';
    RD8_stg  := '0';
    RD9_stg  := '0';
    RD10_stg := '0';
    RD11_stg := '0';
    RD12_stg := '0';
    RD13_stg := '0';
    RD14_stg := '0';
    RD15_stg := '0';
    RD16_stg := '0';
    RD17_stg := '0';
 
  else -- RESET deasserted

    ------------------------------------------------------------
    -- # Synchronization Section                              --
    ------------------------------------------------------------

    if (rising_edge(WCLK_ipd)) then
      -- Synchronizer needs two WCLKs to generate full flag
      RADDR_P2 := RADDR_P1;
      RADDR_P1 := RADDR;
      RADDR_wrap_P2 := RADDR_wrap_P1;
      RADDR_wrap_P1 := not RADDR_wrap;
    end if;

     if (rising_edge(RCLK_ipd)) then
      -- Synchronizer needs two RCLKs to generate empty flag
      WADDR_P2 := WADDR_P1;
      WADDR_P1 := WADDR;
      WADDR_wrap_P2 := WADDR_wrap_P1;
      WADDR_wrap_P1 := WADDR_wrap;
    end if;

    ------------------------------------------------------------
    -- # Write Functional Section                             --
    ------------------------------------------------------------

    if (TO_X01(WCLK_ipd) = 'X' and (WCLK_ipd'event or RESET_ipd'event)) then
--      if (TO_X01(WCLK_previous) /= 'X' or
      if (WCLK_ipd'last_active = now or
          TO_X01(WCLK_ipd'last_value) /= 'X') then
        assert false
          report "WCLK went unknown"
          severity Warning;
      end if;
    elsif (rising_edge(WCLK_ipd)) then
      if ((TO_X01(WBLK_ipd) = '0') and (TO_X01(WEN_ipd) = '0')) then
        if (FULL_zd = '0' or (FULL_zd = '1' and FSTOP_delayed = '0')) then
          case (wwidth) is 
            when 1 =>
              MEM_TMP(WADDR) := WD0_delayed;
              increment_address_counter(WADDR, WADDR_wrap, wwidth, FULL_zd, FSTOP_delayed);
            when 2 =>
              MEM_TMP(WADDR * 2 + 0) := WD0_delayed;
              MEM_TMP(WADDR * 2 + 1) := WD1_delayed;
              increment_address_counter(WADDR, WADDR_wrap, wwidth, FULL_zd, FSTOP_delayed);
            when 4 =>
              MEM_TMP(WADDR * 4 + 0) := WD0_delayed;
              MEM_TMP(WADDR * 4 + 1) := WD1_delayed;
              MEM_TMP(WADDR * 4 + 2) := WD2_delayed;
              MEM_TMP(WADDR * 4 + 3) := WD3_delayed;
              increment_address_counter(WADDR, WADDR_wrap, wwidth, FULL_zd, FSTOP_delayed);
            when 9 =>
              MEM_TMP(WADDR * 8 + 0) := WD0_delayed;
              MEM_TMP(WADDR * 8 + 1) := WD1_delayed;
              MEM_TMP(WADDR * 8 + 2) := WD2_delayed;
              MEM_TMP(WADDR * 8 + 3) := WD3_delayed;
              MEM_TMP(WADDR * 8 + 4) := WD4_delayed;
              MEM_TMP(WADDR * 8 + 5) := WD5_delayed;
              MEM_TMP(WADDR * 8 + 6) := WD6_delayed;
              MEM_TMP(WADDR * 8 + 7) := WD7_delayed;
              MEM9_TMP(WADDR) := WD8_delayed;
              increment_address_counter(WADDR, WADDR_wrap, wwidth, FULL_zd, FSTOP_delayed);
            when 18 =>
              MEM_TMP(WADDR * 16 + 0) := WD0_delayed;
              MEM_TMP(WADDR * 16 + 1) := WD1_delayed;
              MEM_TMP(WADDR * 16 + 2) := WD2_delayed;
              MEM_TMP(WADDR * 16 + 3) := WD3_delayed;
              MEM_TMP(WADDR * 16 + 4) := WD4_delayed;
              MEM_TMP(WADDR * 16 + 5) := WD5_delayed;
              MEM_TMP(WADDR * 16 + 6) := WD6_delayed;
              MEM_TMP(WADDR * 16 + 7) := WD7_delayed;
              MEM9_TMP(WADDR*2 +0) := WD8_delayed;
              MEM_TMP(WADDR * 16 + 8) := WD9_delayed;
              MEM_TMP(WADDR * 16 + 9) := WD10_delayed;
              MEM_TMP(WADDR * 16 + 10) := WD11_delayed;
              MEM_TMP(WADDR * 16 + 11) := WD12_delayed;
              MEM_TMP(WADDR * 16 + 12) := WD13_delayed;
              MEM_TMP(WADDR * 16 + 13) := WD14_delayed;
              MEM_TMP(WADDR * 16 + 14) := WD15_delayed;
              MEM_TMP(WADDR * 16 + 15) := WD16_delayed;
              MEM9_TMP(WADDR * 2 + 1) := WD17_delayed;
              increment_address_counter(WADDR, WADDR_wrap, wwidth, FULL_zd, FSTOP_delayed);
            when others =>
              assert false
              report "Invalid Write port width configuration."
                severity Warning;
          end case;

        elsif (FSTOP_ipd = 'X') then
            assert false 
              report "FSTOP is unknown. When FIFO is EMPTY, to stop writing set FSTOP=1 or to overwrite set FSTOP=0"
              severity Warning;
        end if; -- not(FULL and FSTOP)

      else
        if (TO_X01(WBLK_ipd) = 'X' and (TO_X01(WEN_ipd) = '0' or
                                        TO_X01(WEN_ipd) = 'X')) then
          if ((WBLK_ipd'last_active = now or TO_X01(WBLK_ipd'last_value) /= 'X')
              and issue_WBLK = '0') then
            assert false
              report "WBLK signal is unknown."
              severity Warning;
            issue_WBLK := '1';
          end if;
        end if;
        if(TO_X01(WEN_ipd) = 'X' and (TO_X01(WBLK_ipd) = '0' or
                                      TO_X01(WBLK_ipd) = 'X')) then
          if ((WEN_ipd'last_active = now or TO_X01(WEN_ipd'last_value) /= 'X')
              and issue_WEN = '0') then
            assert false
              report "WEN signal is unknown."
              severity Warning;
            issue_WEN := '1';
          end if;
        end if;
      end if;
        fifo_flags(EMPTY_zd, AEMPTY_zd, FULL_zd, AFULL_zd, RADDR, RADDR_P2, 
                 RADDR_wrap, RADDR_wrap_P2, WADDR, WADDR_P2, WADDR_wrap, 
                 WADDR_wrap_P2, afullvalue, aemptyvalue, MAX_depth, wwidth,
                   rwidth, wwidth_bit, rwidth_bit);
        if (afullvalue < 0 and issue_AFVAL = '0') then

          if (TO_X01(AFVAL11_ipd) = 'X') then
            assert false
              report "AFVAL11 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL10_ipd) = 'X') then
            assert false
              report "AFVAL10 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL9_ipd) = 'X') then
            assert false
              report "AFVAL9 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL8_ipd) = 'X') then
            assert false
              report "AFVAL8 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL7_ipd) = 'X') then
            assert false
              report "AFVAL7 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL6_ipd) = 'X') then
            assert false
              report "AFVAL6 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL5_ipd) = 'X') then
            assert false
              report "AFVAL5 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL4_ipd) = 'X') then
            assert false
              report "AFVAL4 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL3_ipd) = 'X') then
            assert false
              report "AFVAL3 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL2_ipd) = 'X') then
            assert false
              report "AFVAL2 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL1_ipd) = 'X') then
            assert false
              report "AFVAL1 is unknown" severity warning;
          end if;
          if (TO_X01(AFVAL0_ipd) = 'X') then
            assert false
              report "AFVAL0 is unknown" severity warning;
          end if;
          assert false
            report "Holding the value of AFULL flag" severity warning;
          issue_AFVAL := '1';
        elsif (afullvalue >= 0) then
          issue_AFVAL := '0'  ;
        end if;
        
    end if; -- Rising WCLK edge

    --------------------------------------------------------------------
    -- # Read Functional Section                                      --
    --------------------------------------------------------------------

    if (TO_X01(RCLK_ipd) = 'X' and (RCLK_ipd'event or RESET_ipd'event or
                                    REN_ipd'event or RBLK_ipd'event)) then
      if (RCLK_ipd'last_active = now or
          TO_X01(RCLK_ipd'last_value) /= 'X') then
        assert false
          report "RCLK went unknown"
          severity Warning;
      end if;
      if ((TO_X01(REN_ipd) = '1') and (TO_X01(RBLK_ipd) = '0')) then
        RD0_zd   := 'X';
        RD1_zd   := 'X';
        RD2_zd   := 'X';
        RD3_zd   := 'X';
        RD4_zd   := 'X';
        RD5_zd   := 'X';
        RD6_zd   := 'X';
        RD7_zd   := 'X';
        RD8_zd   := 'X';
        RD9_zd   := 'X';
        RD10_zd  := 'X';
        RD11_zd  := 'X';
        RD12_zd  := 'X';
        RD13_zd  := 'X';
        RD14_zd  := 'X';
        RD15_zd  := 'X';
        RD16_zd  := 'X';
        RD17_zd  := 'X';
      end if;
      elsif (rising_edge(RCLK_ipd)) then
      -- fifo read data pipelining
      if (TO_X01(RPIPE_delayed) = '1') then -- Pipelining on
        RD0_zd  := RD0_stg;
        RD1_zd  := RD1_stg;
        RD2_zd  := RD2_stg;
        RD3_zd  := RD3_stg;
        RD4_zd  := RD4_stg;
        RD5_zd  := RD5_stg;
        RD6_zd  := RD6_stg;
        RD7_zd  := RD7_stg;
        RD8_zd  := RD8_stg;
        RD9_zd  := RD9_stg;
        RD10_zd := RD10_stg;
        RD11_zd := RD11_stg;
        RD12_zd := RD12_stg;
        RD13_zd := RD13_stg;
        RD14_zd := RD14_stg;
        RD15_zd := RD15_stg;
        RD16_zd := RD16_stg;
        RD17_zd := RD17_stg;
      elsif (TO_X01(RPIPE_delayed) = 'X') then
        assert false
        report "RPIPE signal unknown."
        severity Warning;
        RD0_zd  := 'X';
        RD1_zd  := 'X';
        RD2_zd  := 'X';
        RD3_zd  := 'X';
        RD4_zd  := 'X';
        RD5_zd  := 'X';
        RD6_zd  := 'X';
        RD7_zd  := 'X';
        RD8_zd  := 'X';
        RD9_zd  := 'X';
        RD10_zd := 'X';
        RD11_zd := 'X';
        RD12_zd := 'X';
        RD13_zd := 'X';
        RD14_zd := 'X';
        RD15_zd := 'X';
        RD16_zd := 'X';
        RD17_zd := 'X';
      end if;
      -- fifo read and flag control logic
      if ((TO_X01(REN_ipd) = '1') and (TO_X01(RBLK_ipd) = '0')) then
        if (EMPTY_zd = '0' or (EMPTY_zd = '1' and ESTOP_delayed = '0')) then
          if (TO_X01(RPIPE_delayed) = '0') then -- Pipelining off
            case (rwidth) is
              when 1  =>
                RD0_zd  := MEM_TMP(RADDR);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 2 =>
                RD0_zd  := MEM_TMP(RADDR * 2 + 0);
                RD1_zd  := MEM_TMP(RADDR * 2 + 1);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 4 =>
                RD0_zd  := MEM_TMP(RADDR * 4 + 0);
                RD1_zd  := MEM_TMP(RADDR * 4 + 1);
                RD2_zd  := MEM_TMP(RADDR * 4 + 2);
                RD3_zd  := MEM_TMP(RADDR * 4 + 3);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 9 =>
                RD0_zd  := MEM_TMP(RADDR * 8 + 0);
                RD1_zd  := MEM_TMP(RADDR * 8 + 1);
                RD2_zd  := MEM_TMP(RADDR * 8 + 2);
                RD3_zd  := MEM_TMP(RADDR * 8 + 3);
                RD4_zd  := MEM_TMP(RADDR * 8 + 4);
                RD5_zd  := MEM_TMP(RADDR * 8 + 5);
                RD6_zd  := MEM_TMP(RADDR * 8 + 6);
                RD7_zd  := MEM_TMP(RADDR * 8 + 7);
                RD8_zd  := MEM9_TMP(RADDR);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 18 =>
                RD0_zd  := MEM_TMP(RADDR * 16 + 0);
                RD1_zd  := MEM_TMP(RADDR * 16 + 1);
                RD2_zd  := MEM_TMP(RADDR * 16 + 2);
                RD3_zd  := MEM_TMP(RADDR * 16 + 3);
                RD4_zd  := MEM_TMP(RADDR * 16 + 4);
                RD5_zd  := MEM_TMP(RADDR * 16 + 5);
                RD6_zd  := MEM_TMP(RADDR * 16 + 6);
                RD7_zd  := MEM_TMP(RADDR * 16 + 7);
                RD8_zd  := MEM9_TMP(RADDR*2 +0);
                RD9_zd  := MEM_TMP(RADDR * 16 + 8);
                RD10_zd := MEM_TMP(RADDR * 16 + 9);
                RD11_zd := MEM_TMP(RADDR * 16 + 10);
                RD12_zd := MEM_TMP(RADDR * 16 + 11);
                RD13_zd := MEM_TMP(RADDR * 16 + 12);
                RD14_zd := MEM_TMP(RADDR * 16 + 13);
                RD15_zd := MEM_TMP(RADDR * 16 + 14);
                RD16_zd := MEM_TMP(RADDR * 16 + 15);
                RD17_zd := MEM9_TMP(RADDR * 2 + 1);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when others =>
                assert false
                report "Illegal Read port width configuration"
                severity Warning;
            end case;
          elsif (TO_X01(RPIPE_delayed) = '1') then -- Pipelining on
            case (rwidth) is
              when 1  =>
                RD0_stg  := MEM_TMP(RADDR);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 2 =>
                RD0_stg  := MEM_TMP(RADDR * 2 + 0);
                RD1_stg  := MEM_TMP(RADDR * 2 + 1);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 4 =>
                RD0_stg  := MEM_TMP(RADDR * 4 + 0);
                RD1_stg  := MEM_TMP(RADDR * 4 + 1);
                RD2_stg  := MEM_TMP(RADDR * 4 + 2);
                RD3_stg  := MEM_TMP(RADDR * 4 + 3);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when 9 =>
                RD0_stg  := MEM_TMP(RADDR * 8 + 0);
                RD1_stg  := MEM_TMP(RADDR * 8 + 1);
                RD2_stg  := MEM_TMP(RADDR * 8 + 2);
                RD3_stg  := MEM_TMP(RADDR * 8 + 3);
                RD4_stg  := MEM_TMP(RADDR * 8 + 4);
                RD5_stg  := MEM_TMP(RADDR * 8 + 5);
                RD6_stg  := MEM_TMP(RADDR * 8 + 6);
                RD7_stg  := MEM_TMP(RADDR * 8 + 7);
                RD8_stg  := MEM9_TMP(RADDR);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed); 
              when 18 =>
                RD0_stg  := MEM_TMP(RADDR * 16 + 0);
                RD1_stg  := MEM_TMP(RADDR * 16 + 1);
                RD2_stg  := MEM_TMP(RADDR * 16 + 2);
                RD3_stg  := MEM_TMP(RADDR * 16 + 3);
                RD4_stg  := MEM_TMP(RADDR * 16 + 4);
                RD5_stg  := MEM_TMP(RADDR * 16 + 5);
                RD6_stg  := MEM_TMP(RADDR * 16 + 6);
                RD7_stg  := MEM_TMP(RADDR * 16 + 7);
                RD8_stg  := MEM9_TMP(RADDR*2   + 0);
                RD9_stg  := MEM_TMP(RADDR * 16 + 8);
                RD10_stg := MEM_TMP(RADDR * 16 + 9);
                RD11_stg := MEM_TMP(RADDR * 16 + 10);
                RD12_stg := MEM_TMP(RADDR * 16 + 11);
                RD13_stg := MEM_TMP(RADDR * 16 + 12);
                RD14_stg := MEM_TMP(RADDR * 16 + 13);
                RD15_stg := MEM_TMP(RADDR * 16 + 14);
                RD16_stg := MEM_TMP(RADDR * 16 + 15);
                RD17_stg := MEM9_TMP(RADDR * 2 + 1);
                increment_address_counter(RADDR, RADDR_wrap, rwidth, EMPTY_zd, ESTOP_delayed);
              when others =>
                assert false
                report "Illegal Read port width configuration"
                  severity Warning;
            end case;
          end if; -- Pipelining
        elsif (ESTOP_ipd = 'X') then
            assert false 
              report "ESTOP is unknown. When FIFO is EMPTY, to stop reading set ESTOP=1 or to continue reading old data set ESTOP=0"
              severity warning;
            issue_ESTOP := '1';
        end if; -- EMPTY
      else
        if(TO_X01(RBLK_ipd) = 'X' and (TO_X01(REN_ipd) = '1' or
                                       TO_X01(REN_ipd) = 'X')) then
          if ((RBLK_ipd'last_active = now or TO_X01(RBLK_ipd'last_value) /= 'X')
              and issue_RBLK = '0') then
            assert false
              report "RBLK signal is unknown."
              severity Warning;
            issue_RBLK := '1';
          end if;
        end if;
        if(TO_X01(REN_ipd) = 'X' and (TO_X01(RBLK_ipd) = '0' or
                                      TO_X01(RBLK_ipd) = 'X')) then
          if ((REN_ipd'last_active = now or TO_X01(REN_ipd'last_value) /= 'X')
            and issue_REN = '0') then
            assert false
              report "REN signal is unknown."
              severity Warning;
            issue_REN := '1';
          end if;
        end if;
      end if;
    fifo_flags(EMPTY_zd, AEMPTY_zd, FULL_zd, AFULL_zd, RADDR, RADDR_P2, 
               RADDR_wrap, RADDR_wrap_P2, WADDR, WADDR_P2, WADDR_wrap, 
               WADDR_wrap_P2, afullvalue, aemptyvalue, MAX_depth, wwidth, rwidth, wwidth_bit, rwidth_bit);

    if (aemptyvalue < 0 and issue_AEVAL = '0' ) then
      if (TO_X01(AEVAL11_ipd) = 'X') then
        assert false
          report "AEVAL11 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL10_ipd) = 'X') then
        assert false
          report "AEVAL10 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL9_ipd) = 'X') then
        assert false
          report "AEVAL9 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL8_ipd) = 'X') then
        assert false
          report "AEVAL8 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL7_ipd) = 'X') then
        assert false
          report "AEVAL7 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL6_ipd) = 'X') then
        assert false
          report "AEVAL6 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL5_ipd) = 'X') then
        assert false
          report "AEVAL5 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL4_ipd) = 'X') then
        assert false
          report "AEVAL4 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL3_ipd) = 'X') then
        assert false
          report "AEVAL3 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL2_ipd) = 'X') then
        assert false
          report "AEVAL2 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL1_ipd) = 'X') then
        assert false
          report "AEVAL1 is unknown" severity warning;
      end if;
      if (TO_X01(AEVAL0_ipd) = 'X') then
        assert false
          report "AEVAL0 is unknown" severity warning;
      end if;
          assert false
            report "Holding the value of AEMPTY flag" severity warning;
      issue_AEVAL := '1';
    elsif (aemptyvalue >= 0) then
      issue_AEVAL := '0'  ;
      
    end if;
  end if; -- rising RCLK edge

 end if; -- RESET deasserted

  WD0_delayed  := WD0_ipd;
  WD1_delayed  := WD1_ipd;
  WD2_delayed  := WD2_ipd;
  WD3_delayed  := WD3_ipd;
  WD4_delayed  := WD4_ipd;
  WD5_delayed  := WD5_ipd;
  WD6_delayed  := WD6_ipd;
  WD7_delayed  := WD7_ipd;
  WD8_delayed  := WD8_ipd;
  WD9_delayed  := WD9_ipd;
  WD10_delayed  := WD10_ipd;
  WD11_delayed  := WD11_ipd;
  WD12_delayed  := WD12_ipd;
  WD13_delayed  := WD13_ipd;
  WD14_delayed  := WD14_ipd;
  WD15_delayed  := WD15_ipd;
  WD16_delayed  := WD16_ipd;
  WD17_delayed  := WD17_ipd;
  ESTOP_delayed := ESTOP_ipd;
  FSTOP_delayed := FSTOP_ipd;

  if (WCLK_ipd'event) then
    WCLK_previous := WCLK_ipd;
  end if;

  if (RCLK_ipd'event) then
    RCLK_previous := RCLK_ipd;
  end if;

if(WBLK_ipd'event and TO_X01(WBLK_ipd) = 'X') then
  issue_WBLK := '0';
end if;
if(RBLK_ipd'event and TO_X01(RBLK_ipd) = 'X') then
  issue_RBLK := '0';
end if;
if(WEN_ipd'event and TO_X01(WEN_ipd) = 'X') then
  issue_WEN := '0';
end if;
if(REN_ipd'event and TO_X01(REN_ipd) = 'X') then
  issue_REN := '0';
end if;
if(ESTOP_ipd'event and TO_X01(ESTOP_ipd) = 'X') then
  issue_ESTOP := '0';
end if;
if(FSTOP_ipd'event and TO_X01(FSTOP_ipd) = 'X') then
  issue_FSTOP := '0';
end if;
RPIPE_delayed := RPIPE_ipd;
RESET_delayed := RESET_ipd;

  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

  VitalPathDelay01Z (
    OutSignal     => RD17,
    GlitchData    => RD17_GlitchData,
    OutSignalName => "RD17",
    OutTemp       => RD17_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD17), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD17), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD16,
    GlitchData    => RD16_GlitchData,
    OutSignalName => "RD16",
    OutTemp       => RD16_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD16), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD16), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD15,
    GlitchData    => RD15_GlitchData,
    OutSignalName => "RD15",
    OutTemp       => RD15_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD15), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD15), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );
  
  VitalPathDelay01Z (
    OutSignal     => RD14,
    GlitchData    => RD14_GlitchData,
    OutSignalName => "RD14",
    OutTemp       => RD14_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD14), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD14), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD13,
    GlitchData    => RD13_GlitchData,
    OutSignalName => "RD13",
    OutTemp       => RD13_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD13), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD13), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );
    
  VitalPathDelay01Z (
    OutSignal     => RD12,
    GlitchData    => RD12_GlitchData,
    OutSignalName => "RD12",
    OutTemp       => RD12_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD12), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD12), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD11,
    GlitchData    => RD11_GlitchData,
    OutSignalName => "RD11",
    OutTemp       => RD11_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD11), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD11), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD10,
    GlitchData    => RD10_GlitchData,
    OutSignalName => "RD10",
    OutTemp       => RD10_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD10), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD10), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD9,
    GlitchData    => RD9_GlitchData,
    OutSignalName => "RD9",
    OutTemp       => RD9_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD9), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD9), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD8,
    GlitchData    => RD8_GlitchData,
    OutSignalName => "RD8",
    OutTemp       => RD8_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD8), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD8), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD7,
    GlitchData    => RD7_GlitchData,
    OutSignalName => "RD7",
    OutTemp       => RD7_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD7), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD6,
    GlitchData    => RD6_GlitchData,
    OutSignalName => "RD6",
    OutTemp       => RD6_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD6), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD5,
    GlitchData    => RD5_GlitchData,
    OutSignalName => "RD5",
    OutTemp       => RD5_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD5), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD4,
    GlitchData    => RD4_GlitchData,
    OutSignalName => "RD4",
    OutTemp       => RD4_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD4), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );
  
  VitalPathDelay01Z (
    OutSignal     => RD3,
    GlitchData    => RD3_GlitchData,
    OutSignalName => "RD3",
    OutTemp       => RD3_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD3), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD2,
    GlitchData    => RD2_GlitchData,
    OutSignalName => "RD2",
    OutTemp       => RD2_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD2), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD1,
    GlitchData    => RD1_GlitchData,
    OutSignalName => "RD1",
    OutTemp       => RD1_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD1), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => RD0,
    GlitchData    => RD0_GlitchData,
    OutSignalName => "RD0",
    OutTemp       => RD0_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_RD0), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => EMPTY,
    GlitchData    => EMPTY_GlitchData,
    OutSignalName => "EMPTY",
    OutTemp       => EMPTY_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_EMPTY), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_EMPTY), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );


  VitalPathDelay01Z (
    OutSignal     => AEMPTY,
    GlitchData    => AEMPTY_GlitchData,
    OutSignalName => "AEMPTY",
    OutTemp       => AEMPTY_zd,
    Paths         => (0 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_AEMPTY), ( AEMPTY_zd = '1' ) ),
                      1 => (WCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_WCLK_AEMPTY), ( AEMPTY_zd = '0' ) ),
                      2 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_AEMPTY), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => AFULL,
    GlitchData    => AFULL_GlitchData,
    OutSignalName => "AFULL",
    OutTemp       => AFULL_zd,
    Paths         => (0 => (WCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_WCLK_AFULL), ( AFULL_zd = '1' ) ),
                      1 => (RCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RCLK_AFULL), ( AFULL_zd = '0' ) ),
                      2 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_AFULL), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );


  VitalPathDelay01Z (
    OutSignal     => FULL,
    GlitchData    => FULL_GlitchData,
    OutSignalName => "FULL",
    OutTemp       => FULL_zd,
    Paths         => (0 => (WCLK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_WCLK_FULL), TRUE),
                      1 => (RESET_ipd'last_event,
                            VitalExtendToFillDelay(tpd_RESET_FULL), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );



  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_FIFO4K18_VITAL of FIFO4K18 is
   for VITAL_ACT
   end for;
end CFG_FIFO4K18_VITAL;


---- CELL UFROM ----
library IEEE;
library STD;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_timing.all;
use IEEE.VITAL_primitives.all;


use std.textio.all;
use ieee.std_logic_textio.all;

entity UFROM is
  generic (

        TimingChecksOn: Boolean := True;
        InstancePath  : String  := "*";
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        MEMORYFILE    : String;
        DATA_X        : Integer := 1;
        ACT_PROGFILE      : String  := "";

        tipd_ADDR0    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR1    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR2    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR3    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR4    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR5    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR6    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_CLK      : VitalDelayType01 := ( 0.000 ns, 0.000 ns );

        tpd_CLK_DO7   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO6   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO5   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO4   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO3   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO2   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO1   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO0   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );

        tsetup_ADDR6_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR6_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR5_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR5_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR4_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR4_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR3_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR3_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR2_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR2_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR1_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR1_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR0_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR0_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tpw_CLK_posedge                   : VitalDelayType := 0.000 ns;
        tpw_CLK_negedge                   : VitalDelayType := 0.000 ns

       );

  port (
        DO0   :  out Std_ulogic := 'X';
        DO1   :  out Std_ulogic := 'X';
        DO2   :  out Std_ulogic := 'X';
        DO3   :  out Std_ulogic := 'X';
        DO4   :  out Std_ulogic := 'X';
        DO5   :  out Std_ulogic := 'X';
        DO6   :  out Std_ulogic := 'X';
        DO7   :  out Std_ulogic := 'X';
        ADDR0 :  in  Std_ulogic := 'X';
        ADDR1 :  in  Std_ulogic := 'X';
        ADDR2 :  in  Std_ulogic := 'X';
        ADDR3 :  in  Std_ulogic := 'X';
        ADDR4 :  in  Std_ulogic := 'X';
        ADDR5 :  in  Std_ulogic := 'X';
        ADDR6 :  in  Std_ulogic := 'X';
        CLK   :  in  Std_ulogic := 'X'
       );
 
  ATTRIBUTE VITAL_LEVEL0 OF UFROM : entity IS TRUE ;
end UFROM;

------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of UFROM is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal ADDR0_ipd : Std_ulogic := 'X';
   signal ADDR1_ipd : Std_ulogic := 'X';
   signal ADDR2_ipd : Std_ulogic := 'X';
   signal ADDR3_ipd : Std_ulogic := 'X';
   signal ADDR4_ipd : Std_ulogic := 'X';
   signal ADDR5_ipd : Std_ulogic := 'X';
   signal ADDR6_ipd : Std_ulogic := 'X';
   signal CLK_ipd   : Std_ulogic := 'X';
 
   signal  INIT_MEM : std_logic:= '0';
   type MEM_TYPE is array (127 downto 0) of std_logic_vector (7 downto 0);
   
 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WireDelay: block
   begin --  block WireDelay
     VitalWireDelay ( ADDR0_ipd, ADDR0, VitalExtendToFillDelay ( tipd_ADDR0 ) );
     VitalWireDelay ( ADDR1_ipd, ADDR1, VitalExtendToFillDelay ( tipd_ADDR1 ) );
     VitalWireDelay ( ADDR2_ipd, ADDR2, VitalExtendToFillDelay ( tipd_ADDR2 ) );
     VitalWireDelay ( ADDR3_ipd, ADDR3, VitalExtendToFillDelay ( tipd_ADDR3 ) );
     VitalWireDelay ( ADDR4_ipd, ADDR4, VitalExtendToFillDelay ( tipd_ADDR4 ) );
     VitalWireDelay ( ADDR5_ipd, ADDR5, VitalExtendToFillDelay ( tipd_ADDR5 ) );
     VitalWireDelay ( ADDR6_ipd, ADDR6, VitalExtendToFillDelay ( tipd_ADDR6 ) );
     VitalWireDelay ( CLK_ipd,   CLK,   VitalExtendToFillDelay ( tipd_CLK   ) );
   end block WireDelay;

   ---- INITIALIZE MEMORY  ----

   process
   begin
      INIT_MEM <= '1';
      wait;
   end process;

 
   VITALBehavior : process (INIT_MEM, ADDR0_ipd, ADDR1_ipd, ADDR2_ipd, 
                            ADDR3_ipd, ADDR4_ipd, ADDR5_ipd, ADDR6_ipd, CLK_ipd )

      -- Internal variable declarations

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;

     variable DO0_GlitchData : VitalGlitchDataType;
     variable DO1_GlitchData : VitalGlitchDataType;
     variable DO2_GlitchData : VitalGlitchDataType;
     variable DO3_GlitchData : VitalGlitchDataType;
     variable DO4_GlitchData : VitalGlitchDataType;
     variable DO5_GlitchData : VitalGlitchDataType;
     variable DO6_GlitchData : VitalGlitchDataType;
     variable DO7_GlitchData : VitalGlitchDataType;

     variable ADDR : integer := -1;
     variable ADDR_REG : std_logic_vector ( 6 downto 0 );

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-128, -128, 0, 1, -128, -128, 0, 1, -128);

     variable memory_array : MEM_TYPE := (others => (others => 'X'));
     variable inline    : LINE;
     variable indata    : std_logic_vector(7 downto 0);
     variable resdata   : std_logic_vector(7 downto 0);

     variable i         : integer := 0;
     file     memfile   : text is MEMORYFILE;

     -- Last value variables
     variable ADDR6_previous : std_ulogic := '0';
     variable ADDR5_previous : std_ulogic := '0';
     variable ADDR4_previous : std_ulogic := '0';
     variable ADDR3_previous : std_ulogic := '0';
     variable ADDR2_previous : std_ulogic := '0';
     variable ADDR1_previous : std_ulogic := '0';
     variable ADDR0_previous : std_ulogic := '0';

     -- timing check results
     VARIABLE Tviol_ADDR6_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR5_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR4_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR3_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR2_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR1_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR0_CLK_posedge     : STD_ULOGIC := '0';

     VARIABLE Tmkr_ADDR6_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR5_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR4_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR3_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR2_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR1_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR0_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;


     VARIABLE Pviol_CLK      : STD_ULOGIC := '0';
     VARIABLE PInfo_CLK      : VitalPeriodDataType := VitalPeriodDataInit;

   begin -- process VITALBehavior

   ------------------------
   --  Timing Check Section
   ------------------------

     if( TimingChecksOn ) then

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR6_CLK_posedge,
         TimingData             => Tmkr_ADDR6_CLK_posedge,
         TestSignal             => ADDR6_ipd,
         TestSignalName         => "ADDR6",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR6_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR6_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR6_CLK_posedge_posedge,
         HoldLow                => thold_ADDR6_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR5_CLK_posedge,
         TimingData             => Tmkr_ADDR5_CLK_posedge,
         TestSignal             => ADDR5_ipd,
         TestSignalName         => "ADDR5",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR5_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR5_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR5_CLK_posedge_posedge,
         HoldLow                => thold_ADDR5_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR4_CLK_posedge,
         TimingData             => Tmkr_ADDR4_CLK_posedge,
         TestSignal             => ADDR4_ipd,
         TestSignalName         => "ADDR4",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR4_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR4_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR4_CLK_posedge_posedge,
         HoldLow                => thold_ADDR4_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR3_CLK_posedge,
         TimingData             => Tmkr_ADDR3_CLK_posedge,
         TestSignal             => ADDR3_ipd,
         TestSignalName         => "ADDR3",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR3_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR3_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR3_CLK_posedge_posedge,
         HoldLow                => thold_ADDR3_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR2_CLK_posedge,
         TimingData             => Tmkr_ADDR2_CLK_posedge,
         TestSignal             => ADDR2_ipd,
         TestSignalName         => "ADDR2",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR2_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR2_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR2_CLK_posedge_posedge,
         HoldLow                => thold_ADDR2_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR1_CLK_posedge,
         TimingData             => Tmkr_ADDR1_CLK_posedge,
         TestSignal             => ADDR1_ipd,
         TestSignalName         => "ADDR1",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR1_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR1_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR1_CLK_posedge_posedge,
         HoldLow                => thold_ADDR1_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR0_CLK_posedge,
         TimingData             => Tmkr_ADDR0_CLK_posedge,
         TestSignal             => ADDR0_ipd,
         TestSignalName         => "ADDR0",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR0_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR0_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR0_CLK_posedge_posedge,
         HoldLow                => thold_ADDR0_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalPeriodPulseCheck (
         Violation              => Pviol_CLK,
         PeriodData             => PInfo_CLK,
         TestSignal             => CLK_ipd,
         TestSignalName         => "CLK",
         TestDelay              => 0 ns,
         Period                 => 0 ns,
         PulseWidthHigh         => tpw_CLK_posedge,
         PulseWidthLow          => tpw_CLK_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/UFROM",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

        end if;


     if ( INIT_MEM'event and INIT_MEM = '1' ) then
       while (( i <= 127 ) and ( not endfile(memfile))) loop
         readline(memfile, inline);
         read(inline, indata);
         resdata := indata;
         memory_array(i) := resdata;
         i := i + 1;
       end loop;
     end if;


     -- register input address on rising edge of CLK_ipd

     if ( CLK_ipd'event and TO_X01(CLK_ipd) = '1' ) then
       ADDR_REG := ( ADDR6_ipd & ADDR5_ipd & ADDR4_ipd & ADDR3_ipd & ADDR2_ipd & ADDR1_ipd & ADDR0_ipd );
       --convert the registered address into integer to access UFROM array
       ADDR     := ( ( INT( ADDR_REG(6) ) * 64 ) + ( INT( ADDR_REG(5) ) * 32 ) + ( INT( ADDR_REG(4) ) * 16) + 
                     ( INT( ADDR_REG(3) ) * 8  ) + ( INT( ADDR_REG(2) ) * 4  ) + ( INT( ADDR_REG(1) ) * 2 ) + 
                     ( INT( ADDR_REG(0) ) * 1  ) );
       if (ADDR < 0) then
         if (TO_X01(ADDR_REG(6)) = 'X' and TO_X01(ADDR6_previous) /= 'X') then
           assert false
           report ": ADDR6 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(5)) = 'X' and TO_X01(ADDR5_previous) /= 'X') then
           assert false
           report ": ADDR5 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(4)) = 'X' and TO_X01(ADDR4_previous) /= 'X') then
           assert false
           report ": ADDR4 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(3)) = 'X' and TO_X01(ADDR3_previous) /= 'X') then
           assert false
           report ": ADDR3 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(2)) = 'X' and TO_X01(ADDR2_previous) /= 'X') then
           assert false
           report ": ADDR2 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(1)) = 'X' and TO_X01(ADDR1_previous) /= 'X') then
           assert false
           report ": ADDR1 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(0)) = 'X' and TO_X01(ADDR0_previous) /= 'X') then
           assert false
           report ": ADDR0 went unknown"
           severity Warning;
         end if;
       end if;
       ADDR6_previous := ADDR_REG(6);
       ADDR5_previous := ADDR_REG(5);
       ADDR4_previous := ADDR_REG(4);
       ADDR3_previous := ADDR_REG(3);
       ADDR2_previous := ADDR_REG(2);
       ADDR1_previous := ADDR_REG(1);
       ADDR0_previous := ADDR_REG(0);

       -- users can turn-off data being driven to "X" on posedge CLK_ipd, by setting DATA_X to 0
       if ( DATA_X = 1 ) then
         DO7_zd := 'X';
         DO6_zd := 'X';
         DO5_zd := 'X';
         DO4_zd := 'X';
         DO3_zd := 'X';
         DO2_zd := 'X';
         DO1_zd := 'X';
         DO0_zd := 'X';
       end if;
     end if;


     -- update DO only on falling edge of CLK_ipd    

     if ( CLK_ipd'event and TO_X01(CLK_ipd) = '0' ) then
       if (ADDR < 0) then
         DO7_zd := 'X';
         DO6_zd := 'X';
         DO5_zd := 'X';
         DO4_zd := 'X';
         DO3_zd := 'X';
         DO2_zd := 'X';
         DO1_zd := 'X';
         DO0_zd := 'X';
       else
         DO0_zd := memory_array(ADDR)(0);
         DO1_zd := memory_array(ADDR)(1);
         DO2_zd := memory_array(ADDR)(2);
         DO3_zd := memory_array(ADDR)(3);
         DO4_zd := memory_array(ADDR)(4);
         DO5_zd := memory_array(ADDR)(5);
         DO6_zd := memory_array(ADDR)(6);
         DO7_zd := memory_array(ADDR)(7);
       end if;
     end if;

     -------------------------------------------------------------
     --              Path Delay Section                         --
     -------------------------------------------------------------

     VitalPathDelay01Z (
       OutSignal     => DO0,
       GlitchData    => DO0_GlitchData,
       OutSignalName => "DO0",
       OutTemp       => DO0_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO0), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );
    
     VitalPathDelay01Z (
       OutSignal     => DO1,
       GlitchData    => DO1_GlitchData,
       OutSignalName => "DO1",
       OutTemp       => DO1_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO1), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO2,
       GlitchData    => DO2_GlitchData,
       OutSignalName => "DO2",
       OutTemp       => DO2_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO2), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO3,
       GlitchData    => DO3_GlitchData,
       OutSignalName => "DO3",
       OutTemp       => DO3_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO3), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO4,
       GlitchData    => DO4_GlitchData,
       OutSignalName => "DO4",
       OutTemp       => DO4_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO4), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO5,
       GlitchData    => DO5_GlitchData,
       OutSignalName => "DO5",
       OutTemp       => DO5_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO5), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO6,
       GlitchData    => DO6_GlitchData,
       OutSignalName => "DO6",
       OutTemp       => DO6_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO6), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO7,
       GlitchData    => DO7_GlitchData,
       OutSignalName => "DO7",
       OutTemp       => DO7_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO7), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

   end process VITALBehavior;

end VITAL_ACT;

configuration CFG_UFROM_VITAL of UFROM is
  for VITAL_ACT
  end for;
end CFG_UFROM_VITAL;



---- CELL UFROMH ----
library IEEE;
library STD;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use IEEE.VITAL_timing.all;
use IEEE.VITAL_primitives.all;


use std.textio.all;
use ieee.std_logic_textio.all;

entity UFROMH is
  generic (

        TimingChecksOn: Boolean := True;
        InstancePath  : String  := "*";
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        MEMORYFILE    : String;
        DATA_X        : Integer := 1;
        ACT_PROGFILE      : String  := "";

        tipd_ADDR0    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR1    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR2    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR3    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR4    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR5    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_ADDR6    : VitalDelayType01 := ( 0.000 ns, 0.000 ns );
        tipd_CLK      : VitalDelayType01 := ( 0.000 ns, 0.000 ns );

        tpd_CLK_DO7   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO6   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO5   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO4   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO3   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO2   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO1   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );
        tpd_CLK_DO0   : VitalDelayType01 := ( 0.100 ns, 0.100 ns );

        tsetup_ADDR6_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR6_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR6_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR5_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR5_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR5_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR4_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR4_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR4_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR3_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR3_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR3_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR2_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR2_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR2_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR1_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR1_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR1_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tsetup_ADDR0_CLK_posedge_posedge  : VitalDelayType := 0.000 ns;
        tsetup_ADDR0_CLK_negedge_posedge  : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_posedge_posedge   : VitalDelayType := 0.000 ns;
        thold_ADDR0_CLK_negedge_posedge   : VitalDelayType := 0.000 ns;

        tpw_CLK_posedge                   : VitalDelayType := 0.000 ns;
        tpw_CLK_negedge                   : VitalDelayType := 0.000 ns

       );

  port (
        DO0   :  out Std_ulogic := 'X';
        DO1   :  out Std_ulogic := 'X';
        DO2   :  out Std_ulogic := 'X';
        DO3   :  out Std_ulogic := 'X';
        DO4   :  out Std_ulogic := 'X';
        DO5   :  out Std_ulogic := 'X';
        DO6   :  out Std_ulogic := 'X';
        DO7   :  out Std_ulogic := 'X';
        ADDR0 :  in  Std_ulogic := 'X';
        ADDR1 :  in  Std_ulogic := 'X';
        ADDR2 :  in  Std_ulogic := 'X';
        ADDR3 :  in  Std_ulogic := 'X';
        ADDR4 :  in  Std_ulogic := 'X';
        ADDR5 :  in  Std_ulogic := 'X';
        ADDR6 :  in  Std_ulogic := 'X';
        CLK   :  in  Std_ulogic := 'X'
       );
 
  ATTRIBUTE VITAL_LEVEL0 OF UFROMH : entity IS TRUE ;
end UFROMH;

------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of UFROMH is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal ADDR0_ipd : Std_ulogic := 'X';
   signal ADDR1_ipd : Std_ulogic := 'X';
   signal ADDR2_ipd : Std_ulogic := 'X';
   signal ADDR3_ipd : Std_ulogic := 'X';
   signal ADDR4_ipd : Std_ulogic := 'X';
   signal ADDR5_ipd : Std_ulogic := 'X';
   signal ADDR6_ipd : Std_ulogic := 'X';
   signal CLK_ipd   : Std_ulogic := 'X';
 
   signal  INIT_MEM : std_logic:= '0';
   type MEM_TYPE is array (127 downto 0) of std_logic_vector (7 downto 0);
   
 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WireDelay: block
   begin --  block WireDelay
     VitalWireDelay ( ADDR0_ipd, ADDR0, VitalExtendToFillDelay ( tipd_ADDR0 ) );
     VitalWireDelay ( ADDR1_ipd, ADDR1, VitalExtendToFillDelay ( tipd_ADDR1 ) );
     VitalWireDelay ( ADDR2_ipd, ADDR2, VitalExtendToFillDelay ( tipd_ADDR2 ) );
     VitalWireDelay ( ADDR3_ipd, ADDR3, VitalExtendToFillDelay ( tipd_ADDR3 ) );
     VitalWireDelay ( ADDR4_ipd, ADDR4, VitalExtendToFillDelay ( tipd_ADDR4 ) );
     VitalWireDelay ( ADDR5_ipd, ADDR5, VitalExtendToFillDelay ( tipd_ADDR5 ) );
     VitalWireDelay ( ADDR6_ipd, ADDR6, VitalExtendToFillDelay ( tipd_ADDR6 ) );
     VitalWireDelay ( CLK_ipd,   CLK,   VitalExtendToFillDelay ( tipd_CLK   ) );
   end block WireDelay;

   ---- INITIALIZE MEMORY  ----

   process
   begin
      INIT_MEM <= '1';
      wait;
   end process;

 
   VITALBehavior : process (INIT_MEM, ADDR0_ipd, ADDR1_ipd, ADDR2_ipd, 
                            ADDR3_ipd, ADDR4_ipd, ADDR5_ipd, ADDR6_ipd, CLK_ipd )

      -- Internal variable declarations

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;

     variable DO0_GlitchData : VitalGlitchDataType;
     variable DO1_GlitchData : VitalGlitchDataType;
     variable DO2_GlitchData : VitalGlitchDataType;
     variable DO3_GlitchData : VitalGlitchDataType;
     variable DO4_GlitchData : VitalGlitchDataType;
     variable DO5_GlitchData : VitalGlitchDataType;
     variable DO6_GlitchData : VitalGlitchDataType;
     variable DO7_GlitchData : VitalGlitchDataType;

     variable ADDR : integer := -1;
     variable ADDR_REG : std_logic_vector ( 6 downto 0 );

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT : SL_TO_INT := (-128, -128, 0, 1, -128, -128, 0, 1, -128);

     variable memory_array : MEM_TYPE := (others => (others => 'X'));
     variable inline    : LINE;
     variable indata    : std_logic_vector(7 downto 0);
     variable resdata   : std_logic_vector(7 downto 0);

     variable i         : integer := 0;
     file     memfile   : text is MEMORYFILE;

     -- Last value variables
     variable ADDR6_previous : std_ulogic := '0';
     variable ADDR5_previous : std_ulogic := '0';
     variable ADDR4_previous : std_ulogic := '0';
     variable ADDR3_previous : std_ulogic := '0';
     variable ADDR2_previous : std_ulogic := '0';
     variable ADDR1_previous : std_ulogic := '0';
     variable ADDR0_previous : std_ulogic := '0';

     -- timing check results
     VARIABLE Tviol_ADDR6_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR5_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR4_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR3_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR2_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR1_CLK_posedge     : STD_ULOGIC := '0';
     VARIABLE Tviol_ADDR0_CLK_posedge     : STD_ULOGIC := '0';

     VARIABLE Tmkr_ADDR6_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR5_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR4_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR3_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR2_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR1_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;
     VARIABLE Tmkr_ADDR0_CLK_posedge      : VitalTimingDataType := VitalTimingDataInit;


     VARIABLE Pviol_CLK      : STD_ULOGIC := '0';
     VARIABLE PInfo_CLK      : VitalPeriodDataType := VitalPeriodDataInit;

   begin -- process VITALBehavior

   ------------------------
   --  Timing Check Section
   ------------------------

     if( TimingChecksOn ) then

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR6_CLK_posedge,
         TimingData             => Tmkr_ADDR6_CLK_posedge,
         TestSignal             => ADDR6_ipd,
         TestSignalName         => "ADDR6",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR6_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR6_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR6_CLK_posedge_posedge,
         HoldLow                => thold_ADDR6_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR5_CLK_posedge,
         TimingData             => Tmkr_ADDR5_CLK_posedge,
         TestSignal             => ADDR5_ipd,
         TestSignalName         => "ADDR5",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR5_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR5_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR5_CLK_posedge_posedge,
         HoldLow                => thold_ADDR5_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR4_CLK_posedge,
         TimingData             => Tmkr_ADDR4_CLK_posedge,
         TestSignal             => ADDR4_ipd,
         TestSignalName         => "ADDR4",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR4_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR4_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR4_CLK_posedge_posedge,
         HoldLow                => thold_ADDR4_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR3_CLK_posedge,
         TimingData             => Tmkr_ADDR3_CLK_posedge,
         TestSignal             => ADDR3_ipd,
         TestSignalName         => "ADDR3",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR3_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR3_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR3_CLK_posedge_posedge,
         HoldLow                => thold_ADDR3_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR2_CLK_posedge,
         TimingData             => Tmkr_ADDR2_CLK_posedge,
         TestSignal             => ADDR2_ipd,
         TestSignalName         => "ADDR2",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR2_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR2_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR2_CLK_posedge_posedge,
         HoldLow                => thold_ADDR2_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR1_CLK_posedge,
         TimingData             => Tmkr_ADDR1_CLK_posedge,
         TestSignal             => ADDR1_ipd,
         TestSignalName         => "ADDR1",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR1_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR1_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR1_CLK_posedge_posedge,
         HoldLow                => thold_ADDR1_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalSetupHoldCheck (
         Violation              => Tviol_ADDR0_CLK_posedge,
         TimingData             => Tmkr_ADDR0_CLK_posedge,
         TestSignal             => ADDR0_ipd,
         TestSignalName         => "ADDR0",
         TestDelay              => 0 ns,
         RefSignal              => CLK_ipd,
         RefSignalName          => "CLK",
         RefDelay               => 0 ns,
         SetupHigh              => tsetup_ADDR0_CLK_posedge_posedge,
         SetupLow               => tsetup_ADDR0_CLK_negedge_posedge,
         HoldHigh               => thold_ADDR0_CLK_posedge_posedge,
         HoldLow                => thold_ADDR0_CLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => 'R',
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

       VitalPeriodPulseCheck (
         Violation              => Pviol_CLK,
         PeriodData             => PInfo_CLK,
         TestSignal             => CLK_ipd,
         TestSignalName         => "CLK",
         TestDelay              => 0 ns,
         Period                 => 0 ns,
         PulseWidthHigh         => tpw_CLK_posedge,
         PulseWidthLow          => tpw_CLK_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/UFROMH",
         Xon            => Xon,
         MsgOn          => MsgOn,
         MsgSeverity    => WARNING);

        end if;


     if ( INIT_MEM'event and INIT_MEM = '1' ) then
       while (( i <= 127 ) and ( not endfile(memfile))) loop
         readline(memfile, inline);
         read(inline, indata);
         resdata := indata;
         memory_array(i) := resdata;
         i := i + 1;
       end loop;
     end if;


     -- register input address on rising edge of CLK_ipd

     if ( CLK_ipd'event and TO_X01(CLK_ipd) = '1' ) then
       ADDR_REG := ( ADDR6_ipd & ADDR5_ipd & ADDR4_ipd & ADDR3_ipd & ADDR2_ipd & ADDR1_ipd & ADDR0_ipd );
       --convert the registered address into integer to access UFROM array
       ADDR     := ( ( INT( ADDR_REG(6) ) * 64 ) + ( INT( ADDR_REG(5) ) * 32 ) + ( INT( ADDR_REG(4) ) * 16) + 
                     ( INT( ADDR_REG(3) ) * 8  ) + ( INT( ADDR_REG(2) ) * 4  ) + ( INT( ADDR_REG(1) ) * 2 ) + 
                     ( INT( ADDR_REG(0) ) * 1  ) );
       if (ADDR < 0) then
         if (TO_X01(ADDR_REG(6)) = 'X' and TO_X01(ADDR6_previous) /= 'X') then
           assert false
           report ": ADDR6 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(5)) = 'X' and TO_X01(ADDR5_previous) /= 'X') then
           assert false
           report ": ADDR5 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(4)) = 'X' and TO_X01(ADDR4_previous) /= 'X') then
           assert false
           report ": ADDR4 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(3)) = 'X' and TO_X01(ADDR3_previous) /= 'X') then
           assert false
           report ": ADDR3 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(2)) = 'X' and TO_X01(ADDR2_previous) /= 'X') then
           assert false
           report ": ADDR2 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(1)) = 'X' and TO_X01(ADDR1_previous) /= 'X') then
           assert false
           report ": ADDR1 went unknown"
           severity Warning;
         end if;
         if (TO_X01(ADDR_REG(0)) = 'X' and TO_X01(ADDR0_previous) /= 'X') then
           assert false
           report ": ADDR0 went unknown"
           severity Warning;
         end if;
       end if;
       ADDR6_previous := ADDR_REG(6);
       ADDR5_previous := ADDR_REG(5);
       ADDR4_previous := ADDR_REG(4);
       ADDR3_previous := ADDR_REG(3);
       ADDR2_previous := ADDR_REG(2);
       ADDR1_previous := ADDR_REG(1);
       ADDR0_previous := ADDR_REG(0);

       -- users can turn-off data being driven to "X" on posedge CLK_ipd, by setting DATA_X to 0
       if ( DATA_X = 1 ) then
         DO7_zd := 'X';
         DO6_zd := 'X';
         DO5_zd := 'X';
         DO4_zd := 'X';
         DO3_zd := 'X';
         DO2_zd := 'X';
         DO1_zd := 'X';
         DO0_zd := 'X';
       end if;
     end if;


     -- update DO only on falling edge of CLK_ipd    

     if ( CLK_ipd'event and TO_X01(CLK_ipd) = '0' ) then
       if (ADDR < 0) then
         DO7_zd := 'X';
         DO6_zd := 'X';
         DO5_zd := 'X';
         DO4_zd := 'X';
         DO3_zd := 'X';
         DO2_zd := 'X';
         DO1_zd := 'X';
         DO0_zd := 'X';
       else
         DO0_zd := memory_array(ADDR)(0);
         DO1_zd := memory_array(ADDR)(1);
         DO2_zd := memory_array(ADDR)(2);
         DO3_zd := memory_array(ADDR)(3);
         DO4_zd := memory_array(ADDR)(4);
         DO5_zd := memory_array(ADDR)(5);
         DO6_zd := memory_array(ADDR)(6);
         DO7_zd := memory_array(ADDR)(7);
       end if;
     end if;

     -------------------------------------------------------------
     --              Path Delay Section                         --
     -------------------------------------------------------------

     VitalPathDelay01Z (
       OutSignal     => DO0,
       GlitchData    => DO0_GlitchData,
       OutSignalName => "DO0",
       OutTemp       => DO0_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO0), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );
    
     VitalPathDelay01Z (
       OutSignal     => DO1,
       GlitchData    => DO1_GlitchData,
       OutSignalName => "DO1",
       OutTemp       => DO1_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO1), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO2,
       GlitchData    => DO2_GlitchData,
       OutSignalName => "DO2",
       OutTemp       => DO2_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO2), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO3,
       GlitchData    => DO3_GlitchData,
       OutSignalName => "DO3",
       OutTemp       => DO3_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO3), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO4,
       GlitchData    => DO4_GlitchData,
       OutSignalName => "DO4",
       OutTemp       => DO4_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO4), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO5,
       GlitchData    => DO5_GlitchData,
       OutSignalName => "DO5",
       OutTemp       => DO5_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO5), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO6,
       GlitchData    => DO6_GlitchData,
       OutSignalName => "DO6",
       OutTemp       => DO6_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO6), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

     VitalPathDelay01Z (
       OutSignal     => DO7,
       GlitchData    => DO7_GlitchData,
       OutSignalName => "DO7",
       OutTemp       => DO7_zd,
       Paths         => (0 => (CLK_ipd'last_event,
                               VitalExtendToFillDelay(tpd_CLK_DO7), true)),
       DefaultDelay  => VitalZeroDelay01Z,
       Mode          => VitalTransport,
       Xon           => Xon,
       MsgOn         => MsgOn,
       MsgSeverity   => Warning
      );

   end process VITALBehavior;

end VITAL_ACT;

configuration CFG_UFROMH_VITAL of UFROMH is
  for VITAL_ACT
  end for;
end CFG_UFROMH_VITAL;



----- CELL CLKDIVDLY1 -----


--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
--library IEEE;
--use IEEE.VITAL_Timing.all;

-- entity declaration --
--entity CLKDIVDLY1 is
--   generic(
--        TimingChecksOn: Boolean := True;
--        InstancePath: STRING := "*";
--        Xon: Boolean := False;
--        MsgOn: Boolean := True;
--        tipd_CLK         :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYY4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns );
--        tpd_CLK_Y         :  VitalDelayType01 := (  0.1 ns,0.1 ns ));
--
--     port (
--        CLK         : in    STD_ULOGIC;
--        ODIV0       : in    STD_ULOGIC;
--        ODIV1       : in    STD_ULOGIC;
--        ODIV2       : in    STD_ULOGIC;
--        ODIV3       : in    STD_ULOGIC;
--        ODIV4       : in    STD_ULOGIC;
--        DLYY0       : in    STD_ULOGIC;
--        DLYY1       : in    STD_ULOGIC;
--        DLYY2       : in    STD_ULOGIC;
--        DLYY3       : in    STD_ULOGIC;
--        DLYY4       : in    STD_ULOGIC;
--        DLYGL0       : in    STD_ULOGIC;
--        DLYGL1       : in    STD_ULOGIC;
--        DLYGL2       : in    STD_ULOGIC;
--        DLYGL3       : in    STD_ULOGIC;
--        DLYGL4       : in    STD_ULOGIC;
--        GL           : out   STD_ULOGIC;
--        Y            : out   STD_ULOGIC);
--
--  
--attribute VITAL_LEVEL0 of CLKDIVDLY1 : entity is TRUE;
--end CLKDIVDLY1;
--
---- architecture body --
--library IEEE;
--use IEEE.VITAL_Primitives.all;
--architecture VITAL_ACT of CLKDIVDLY1 is
-- attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;
--
--
-- SIGNAL   CLK_ipd          :   STD_ULOGIC;
-- SIGNAL   ODIV0_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV1_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV2_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV3_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV4_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYY0_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYY1_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYY2_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYY3_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYY4_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL0_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL1_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL2_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL3_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL4_ipd        :   STD_ULOGIC;
--
-- SIGNAL DIV           : Integer := 1; -- Divide by a divisor - range 1 to 128
-- SIGNAL YDELAY       : Time := 0.000 ns; -- Additional Global B Delay
-- SIGNAL GLDELAY       : Time := 0.000 ns; -- Additional Global B Delay
-- SIGNAL DIVout        :   STD_ULOGIC;
--
--begin
--  ---------------------
--   --  INPUT PATH DELAYs
--   ---------------------
--   WireDelay : block
--
--   begin
--
--     VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
--     VitalWireDelay (ODIV0_ipd, ODIV0, tipd_ODIV0);
--     VitalWireDelay (ODIV1_ipd, ODIV1, tipd_ODIV1);
--     VitalWireDelay (ODIV2_ipd, ODIV2, tipd_ODIV2);
--     VitalWireDelay (ODIV3_ipd, ODIV3, tipd_ODIV3);
--     VitalWireDelay (ODIV4_ipd, ODIV4, tipd_ODIV4);
--     VitalWireDelay (DLYY0_ipd, DLYY0, tipd_DLYY0);
--     VitalWireDelay (DLYY1_ipd, DLYY1, tipd_DLYY1);
--     VitalWireDelay (DLYY2_ipd, DLYY2, tipd_DLYY2);
--     VitalWireDelay (DLYY3_ipd, DLYY3, tipd_DLYY3);
--     VitalWireDelay (DLYY4_ipd, DLYY4, tipd_DLYY4);
--     VitalWireDelay (DLYGL0_ipd, DLYGL0, tipd_DLYGL0);
--     VitalWireDelay (DLYGL1_ipd, DLYGL1, tipd_DLYGL1);
--     VitalWireDelay (DLYGL2_ipd, DLYGL2, tipd_DLYGL2);
--     VitalWireDelay (DLYGL3_ipd, DLYGL3, tipd_DLYGL3);
--     VitalWireDelay (DLYGL4_ipd, DLYGL4, tipd_DLYGL4);
--
--   end block WireDelay;
--
--  -- #########################################################
--  -- # Behavior Section
--  -- #########################################################
--
----
--  -- Get GL Delay
--  --
--
-- GetGLDelay : process ( DLYGL0_ipd, DLYGL1_ipd, DLYGL2_ipd, DLYGL3_ipd, DLYGL4_ipd)
--   variable DLYGL : STD_ULOGIC_VECTOR(4 downto 0);
--
--  begin
--
--   DLYGL := DLYGL4_ipd & DLYGL3_ipd & DLYGL2_ipd & DLYGL1_ipd & DLYGL0_ipd;
--
--   case DLYGL is
--         when "00000" =>  GLDELAY <= 0.400 ns;
--         when "00001" =>  GLDELAY <= 0.525 ns;
--         when "00010" =>  GLDELAY <= 0.650 ns;
--         when "00011" =>  GLDELAY <= 0.775 ns;
--         when "00100" =>  GLDELAY <= 0.900 ns;
--         when "00101" =>  GLDELAY <= 1.025 ns;
--         when "00110" =>  GLDELAY <= 1.150 ns;
--         when "00111" =>  GLDELAY <= 1.275 ns;
--         when "01000" =>  GLDELAY <= 1.400 ns;
--         when "01001" =>  GLDELAY <= 1.525 ns;
--         when "01010" =>  GLDELAY <= 1.650 ns;
--         when "01011" =>  GLDELAY <= 1.775 ns;
--         when "01100" =>  GLDELAY <= 1.900 ns;
--         when "01101" =>  GLDELAY <= 2.025 ns;
--         when "01110" =>  GLDELAY <= 2.150 ns;
--         when "01111" =>  GLDELAY <= 2.275 ns;
--         when "10000" =>  GLDELAY <= 2.400 ns;
--         when "10001" =>  GLDELAY <= 2.525 ns;
--         when "10010" =>  GLDELAY <= 2.650 ns;
--         when "10011" =>  GLDELAY <= 2.775 ns;
--         when "10100" =>  GLDELAY <= 2.900 ns;
--         when "10101" =>  GLDELAY <= 3.025 ns;
--         when "10110" =>  GLDELAY <= 3.150 ns;
--         when "10111" =>  GLDELAY <= 3.275 ns;
--         when "11000" =>  GLDELAY <= 3.400 ns;
--         when "11001" =>  GLDELAY <= 3.525 ns;
--         when "11010" =>  GLDELAY <= 3.650 ns;
--         when "11011" =>  GLDELAY <= 3.775 ns;
--         when "11100" =>  GLDELAY <= 3.900 ns;
--         when "11101" =>  GLDELAY <= 4.025 ns;
--         when "11110" =>  GLDELAY <= 4.150 ns;
--         when "11111" =>  GLDELAY <= 4.275 ns;
--         when others =>  GLDELAY <= 0.00 ns;
--
--    end case;
--
--  end process GetGLDelay;
--
--  --
--  -- Get YB Delay
--  --
--
-- GetYDelay : process ( DLYY0_ipd, DLYY1_ipd, DLYY2_ipd, DLYY3_ipd, DLYY4_ipd)
--   variable DLYY : STD_ULOGIC_VECTOR(4 downto 0);
--
--  begin
--
--   DLYY := DLYY4_ipd & DLYY3_ipd & DLYY2_ipd & DLYY1_ipd & DLYY0_ipd;
--   case DLYY is
--         when "00000" =>  YDELAY <= 0.400 ns;
--         when "00001" =>  YDELAY <= 0.525 ns;
--         when "00010" =>  YDELAY <= 0.650 ns;
--         when "00011" =>  YDELAY <= 0.775 ns;
--         when "00100" =>  YDELAY <= 0.900 ns;
--         when "00101" =>  YDELAY <= 1.025 ns;
--         when "00110" =>  YDELAY <= 1.150 ns;
--         when "00111" =>  YDELAY <= 1.275 ns;
--         when "01000" =>  YDELAY <= 1.400 ns;
--         when "01001" =>  YDELAY <= 1.525 ns;
--         when "01010" =>  YDELAY <= 1.650 ns;
--         when "01011" =>  YDELAY <= 1.775 ns;
--         when "01100" =>  YDELAY <= 1.900 ns;
--         when "01101" =>  YDELAY <= 2.025 ns;
--         when "01110" =>  YDELAY <= 2.150 ns;
--         when "01111" =>  YDELAY <= 2.275 ns;
--         when "10000" =>  YDELAY <= 2.400 ns;
--         when "10001" =>  YDELAY <= 2.525 ns;
--         when "10010" =>  YDELAY <= 2.650 ns;
--         when "10011" =>  YDELAY <= 2.775 ns;
--         when "10100" =>  YDELAY <= 2.900 ns;
--         when "10101" =>  YDELAY <= 3.025 ns;
--         when "10110" =>  YDELAY <= 3.150 ns;
--         when "10111" =>  YDELAY <= 3.275 ns;
--         when "11000" =>  YDELAY <= 3.400 ns;
--         when "11001" =>  YDELAY <= 3.525 ns;
--         when "11010" =>  YDELAY <= 3.650 ns;
--         when "11011" =>  YDELAY <= 3.775 ns;
--         when "11100" =>  YDELAY <= 3.900 ns;
--         when "11101" =>  YDELAY <= 4.025 ns;
--         when "11110" =>  YDELAY <= 4.150 ns;
--         when "11111" =>  YDELAY <= 4.275 ns;
--         when others =>   YDELAY <= 0.00 ns;
--
--    end case;
--
--end process GetYDelay;
--
--
--   --
--  -- Get DIV value
--  --
--
--  GetDiv : process ( ODIV4_ipd,ODIV3_ipd,ODIV2_ipd,ODIV1_ipd,ODIV0_ipd)
--    variable ODIV  : STD_ULOGIC_VECTOR(4 downto 0);
--    variable DivVal : Integer := 0;
--
--  begin
--    ODIV := ODIV4_ipd&ODIV3_ipd&ODIV2_ipd&ODIV1_ipd&ODIV0_ipd;
--    DivVal := 0;
--    for i in 0 to 4 loop
--      if (ODIV(i) = '1') then
--        DivVal := DivVal + (2**i);
--      end if;
--    end loop;
--
--    DIV <= DivVal + 1;
--
--  end process GetDiv;
--
--
--
--  --
--  --  Output of Divider
--  --  Assumes input 50/50 duty cycle
--  --
--
--  OutDiv : process (CLK_ipd, DIV)
--
--    variable Q         : STD_LOGIC := '0';
--    variable num_edges : Integer   :=  -1;
--
--  begin
--
--
--   if(CLK_ipd'event ) then
--      num_edges := num_edges + 1;
--   end if;
--
--   if(DIV'event) then
--      num_edges := -1;
--   end if;
-- 
--  if( DIV /=1 ) then
--   if (num_edges mod DIV = 1) then
--       Q := not Q;
--   else
--       Q := Q;
--   end if;
--
--  else
--      Q := CLK_ipd;
--  end if;
--
--  DIVout <= Q;
--
-- end process OutDiv;
--
--
--
----
---- get Y output
----
--
-- getY : process(DIVout, YDELAY)
-- begin
--       Y <= DIVout after YDELAY;
-- end process getY;
--
--
----
----  get the GL output value
----
--
--getGL : process(DIVout, GLDELAY)
--
--begin
--
--     GL <= DIVout after GLDELAY;
--
-- end process getGL;
--
--
--end VITAL_ACT;
--
--configuration CFG_CLKDIVDLY1_VITAL of CLKDIVDLY1 is
--   for VITAL_ACT
--   end for;
--end CFG_CLKDIVDLY1_VITAL;
--
------- CELL CLKDIVDLY -----
--
--library IEEE;
--use IEEE.STD_LOGIC_1164.all;
--library IEEE;
--use IEEE.VITAL_Timing.all;
--
---- entity declaration --
--entity CLKDIVDLY is
--   generic(
--        TimingChecksOn: Boolean := True;
--        InstancePath: STRING := "*";
--        Xon: Boolean := False;
--        MsgOn: Boolean := True;
--        tipd_CLK         :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_ODIV4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
--        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns ));
--
--     port (
--        CLK         : in    STD_ULOGIC;
--        ODIV0       : in    STD_ULOGIC;
--        ODIV1       : in    STD_ULOGIC;
--        ODIV2       : in    STD_ULOGIC;
--        ODIV3       : in    STD_ULOGIC;
--        ODIV4       : in    STD_ULOGIC;
--        DLYGL0       : in    STD_ULOGIC;
--        DLYGL1       : in    STD_ULOGIC;
--        DLYGL2       : in    STD_ULOGIC;
--        DLYGL3       : in    STD_ULOGIC;
--        DLYGL4       : in    STD_ULOGIC;
--        GL           : out   STD_ULOGIC
--          );
--
-- 
--attribute VITAL_LEVEL0 of CLKDIVDLY : entity is TRUE;
--end CLKDIVDLY;
--
--
--
---- architecture body --
--library IEEE;
--use IEEE.VITAL_Primitives.all;
--architecture VITAL_ACT of CLKDIVDLY is
-- attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;
--
-- SIGNAL   CLK_ipd          :   STD_ULOGIC;
-- SIGNAL   ODIV0_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV1_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV2_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV3_ipd        :   STD_ULOGIC;
-- SIGNAL   ODIV4_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL0_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL1_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL2_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL3_ipd        :   STD_ULOGIC;
-- SIGNAL   DLYGL4_ipd        :   STD_ULOGIC;
--
-- SIGNAL DIV           : Integer := 1; -- Divide by a divisor - range 1 to 128
-- SIGNAL GLDELAY       : Time := 0.000 ns; -- Additional Global B Delay
-- SIGNAL DIVout        :   STD_ULOGIC;
--
--begin
--
--   ---------------------
--   --  INPUT PATH DELAYs
--   ---------------------
--   WireDelay : block
--
--   begin
--
--     VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
--     VitalWireDelay (ODIV0_ipd, ODIV0, tipd_ODIV0);
--     VitalWireDelay (ODIV1_ipd, ODIV1, tipd_ODIV1);
--     VitalWireDelay (ODIV2_ipd, ODIV2, tipd_ODIV2);
--     VitalWireDelay (ODIV3_ipd, ODIV3, tipd_ODIV3);
--     VitalWireDelay (ODIV4_ipd, ODIV4, tipd_ODIV4);
--     VitalWireDelay (DLYGL0_ipd, DLYGL0, tipd_DLYGL0);
--     VitalWireDelay (DLYGL1_ipd, DLYGL1, tipd_DLYGL1);
--     VitalWireDelay (DLYGL2_ipd, DLYGL2, tipd_DLYGL2);
--     VitalWireDelay (DLYGL3_ipd, DLYGL3, tipd_DLYGL3);
--     VitalWireDelay (DLYGL4_ipd, DLYGL4, tipd_DLYGL4);
--
--   end block WireDelay;
--
-- 
--
--  -- #########################################################
--  -- # Behavior Section
--  -- #########################################################
--
--
--  --
--  -- Get GL Delay
--  --
--
-- GetGLDelay : process ( DLYGL0_ipd, DLYGL1_ipd, DLYGL2_ipd, DLYGL3_ipd, DLYGL4_ipd)
--   variable DLYGL : STD_ULOGIC_VECTOR(4 downto 0);
--
--  begin
--
--   DLYGL := DLYGL4_ipd & DLYGL3_ipd & DLYGL2_ipd & DLYGL1_ipd & DLYGL0_ipd;
--
--   case DLYGL is
--
--         when "00000" =>  GLDELAY <= 0.400 ns;
--         when "00001" =>  GLDELAY <= 0.525 ns;
--         when "00010" =>  GLDELAY <= 0.650 ns;
--         when "00011" =>  GLDELAY <= 0.775 ns;
--         when "00100" =>  GLDELAY <= 0.900 ns;
--         when "00101" =>  GLDELAY <= 1.025 ns;
--         when "00110" =>  GLDELAY <= 1.150 ns;
--         when "00111" =>  GLDELAY <= 1.275 ns;
--         when "01000" =>  GLDELAY <= 1.400 ns;
--         when "01001" =>  GLDELAY <= 1.525 ns;
--         when "01010" =>  GLDELAY <= 1.650 ns;
--         when "01011" =>  GLDELAY <= 1.775 ns;
--         when "01100" =>  GLDELAY <= 1.900 ns;
--         when "01101" =>  GLDELAY <= 2.025 ns;
--         when "01110" =>  GLDELAY <= 2.150 ns;
--         when "01111" =>  GLDELAY <= 2.275 ns;
--         when "10000" =>  GLDELAY <= 2.400 ns;
--         when "10001" =>  GLDELAY <= 2.525 ns;
--         when "10010" =>  GLDELAY <= 2.650 ns;
--         when "10011" =>  GLDELAY <= 2.775 ns;
--         when "10100" =>  GLDELAY <= 2.900 ns;
--         when "10101" =>  GLDELAY <= 3.025 ns;
--         when "10110" =>  GLDELAY <= 3.150 ns;
--         when "10111" =>  GLDELAY <= 3.275 ns;
--         when "11000" =>  GLDELAY <= 3.400 ns;
--         when "11001" =>  GLDELAY <= 3.525 ns;
--         when "11010" =>  GLDELAY <= 3.650 ns;
--         when "11011" =>  GLDELAY <= 3.775 ns;
--         when "11100" =>  GLDELAY <= 3.900 ns;
--         when "11101" =>  GLDELAY <= 4.025 ns;
--         when "11110" =>  GLDELAY <= 4.150 ns;
--         when "11111" =>  GLDELAY <= 4.275 ns;
--         when others =>  GLDELAY <= 0.00 ns;
--
--    end case;
--  end process GetGLDelay;
--
--   --
--  -- Get DIV value
--  --
--
--  GetDiv : process ( ODIV4_ipd,ODIV3_ipd,ODIV2_ipd,ODIV1_ipd,ODIV0_ipd)
--    variable ODIV  : STD_ULOGIC_VECTOR(4 downto 0);
--    variable DivVal : Integer := 0;
--
--  begin
--    ODIV := ODIV4_ipd&ODIV3_ipd&ODIV2_ipd&ODIV1_ipd&ODIV0_ipd;
--    DivVal := 0;
--    for i in 0 to 4 loop
--      if (ODIV(i) = '1') then
--        DivVal := DivVal + (2**i);
--      end if;
--    end loop;
--
--    DIV <= DivVal + 1;
--
--  end process GetDiv;
--
--
-- 
--
--  --
--  --  Output of Divider
--  --  Assumes input 50/50 duty cycle
--  --
--
--  OutDiv : process (CLK_ipd, DIV)
--
--    variable Q         : STD_LOGIC := '0';
--    variable num_edges : Integer   :=  -1;
--
--  begin
--
--
--   if(CLK_ipd'event ) then
--      num_edges := num_edges + 1;
--   end if;
--
--   if(DIV'event) then
--      num_edges := -1;
--    end if;
--
--
--  if( DIV /=1 ) then
--   if (num_edges mod DIV = 1) then
--       Q := not Q;
--   else
--       Q := Q;
--   end if;
--
--  else
--      Q := CLK_ipd;
--  end if;
--
--  DIVout <= Q;
--
-- end process OutDiv;
--
--
----
----  get the GL output value
----
--
--getGL : process(DIVout, GLDELAY)
--
--begin
--
--     GL <= DIVout after GLDELAY;
--
-- end process getGL;
--
--
--end VITAL_ACT;
--
--configuration CFG_CLKDIVDLY_VITAL of CLKDIVDLY is
--   for VITAL_ACT
--   end for;
--end CFG_CLKDIVDLY_VITAL;


----- CELL CLKDLY -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
use IEEE.STD_LOGIC_ARITH.all;

-- entity declaration --
 entity CLKDLY is
   generic(
        TimingChecksOn : Boolean := True;
        InstancePath   : STRING  := "*";
        Xon            : Boolean := False;
        MsgOn          : Boolean := True;
        INTRINSIC_DELAY     : Time             := 0.470 ns;
        PROG_INIT_DELAY     : Time             := 1.610 ns;
        PROG_STEP_INCREMENT : Time             := 0.360 ns;
        tipd_CLK          :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns ));

     port (
        CLK          : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL           : out   STD_ULOGIC
          );


attribute VITAL_LEVEL0 of CLKDLY : entity is TRUE;
end CLKDLY;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKDLY is
 attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

 SIGNAL   CLK_ipd           :   STD_ULOGIC;
 SIGNAL   DLYGL0_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL1_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL2_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL3_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL4_ipd        :   STD_ULOGIC;

 SIGNAL   GLDELAY           :   Time := 0.000 ns; -- Additional Global B Delay

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

     VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
     VitalWireDelay (DLYGL0_ipd, DLYGL0, tipd_DLYGL0);
     VitalWireDelay (DLYGL1_ipd, DLYGL1, tipd_DLYGL1);
     VitalWireDelay (DLYGL2_ipd, DLYGL2, tipd_DLYGL2);
     VitalWireDelay (DLYGL3_ipd, DLYGL3, tipd_DLYGL3);
     VitalWireDelay (DLYGL4_ipd, DLYGL4, tipd_DLYGL4);

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################


  --
  -- Get GL Delay
  --

 GetGLDelay : process ( DLYGL0_ipd, DLYGL1_ipd, DLYGL2_ipd, DLYGL3_ipd, DLYGL4_ipd)
   variable DLYGL : STD_ULOGIC_VECTOR(4 downto 0);
   variable step : integer;
  begin
    DLYGL := DLYGL4_ipd & DLYGL3_ipd & DLYGL2_ipd & DLYGL1_ipd & DLYGL0_ipd;
    if ( IS_X( DLYGL ) ) then
      GLDELAY <= 0.0 ns;
    else
      step := CONV_INTEGER( unsigned( DLYGL ) );
      if ( step = 0 ) then
        GLDELAY <= INTRINSIC_DELAY;
      else
        GLDELAY <= INTRINSIC_DELAY + ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
      end if;
    end if;
  end process GetGLDelay;

--
--  get the GL output value
--

getGL : process(CLK_ipd, GLDELAY)

begin

     GL <= transport CLK_ipd after GLDELAY;

 end process getGL;


end VITAL_ACT;

configuration CFG_CLKDLY_VITAL of CLKDLY is
   for VITAL_ACT
   end for;
end CFG_CLKDLY_VITAL;


----- CELL CLKDLYINT -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
 entity CLKDLYINT is
   generic(
        TimingChecksOn : Boolean := True;
        InstancePath   : STRING  := "*";
        Xon            : Boolean := False;
        MsgOn          : Boolean := True;
        tipd_CLK          :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns ));

     port (
        CLK          : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL           : out   STD_ULOGIC
          );


attribute VITAL_LEVEL0 of CLKDLYINT : entity is TRUE;
end CLKDLYINT;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKDLYINT is
 attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

 SIGNAL   CLK_ipd           :   STD_ULOGIC;
 SIGNAL   CLK_prev          :   STD_ULOGIC;
 SIGNAL   DLYGL0_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL1_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL2_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL3_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL4_ipd        :   STD_ULOGIC;

 SIGNAL   GLDELAY           :   Time := 0.921 ns; -- Additional Global B Delay

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

     VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
     VitalWireDelay (DLYGL0_ipd, DLYGL0, tipd_DLYGL0);
     VitalWireDelay (DLYGL1_ipd, DLYGL1, tipd_DLYGL1);
     VitalWireDelay (DLYGL2_ipd, DLYGL2, tipd_DLYGL2);
     VitalWireDelay (DLYGL3_ipd, DLYGL3, tipd_DLYGL3);
     VitalWireDelay (DLYGL4_ipd, DLYGL4, tipd_DLYGL4);

   end block WireDelay;


  -- #########################################################
  -- # Behavior Section
  -- #########################################################


  --
  --  get the GL output value
  --

  getGL : process(CLK_ipd, GLDELAY)

  begin

     if ( tpd_CLK_GL = VitalZeroDelay01 ) then
       GL <= transport CLK_ipd after GLDELAY;
     else
       GL <= transport CLK_ipd after VitalCalcDelay ( CLK_ipd, CLK_prev, tpd_CLK_GL );
     end if;

     CLK_prev <= CLK_ipd;

  end process getGL;

 end VITAL_ACT;

configuration CFG_CLKDLYINT_VITAL of CLKDLYINT is
   for VITAL_ACT
   end for;
end CFG_CLKDLYINT_VITAL;


----- CELL CLKDLYIO -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
 entity CLKDLYIO is
   generic(
        TimingChecksOn : Boolean := True;
        InstancePath   : STRING  := "*";
        Xon            : Boolean := False;
        MsgOn          : Boolean := True;
        tipd_CLK          :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL0       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL1       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL2       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL3       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tipd_DLYGL4       :  VitalDelayType01 := (  0.0 ns,0.0 ns );
        tpd_CLK_GL        :  VitalDelayType01 := (  0.1 ns,0.1 ns ));

     port (
        CLK          : in    STD_ULOGIC;
        DLYGL0       : in    STD_ULOGIC;
        DLYGL1       : in    STD_ULOGIC;
        DLYGL2       : in    STD_ULOGIC;
        DLYGL3       : in    STD_ULOGIC;
        DLYGL4       : in    STD_ULOGIC;
        GL           : out   STD_ULOGIC
          );


attribute VITAL_LEVEL0 of CLKDLYIO : entity is TRUE;
end CLKDLYIO;


-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CLKDLYIO is
 attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

 SIGNAL   CLK_ipd           :   STD_ULOGIC;
 SIGNAL   CLK_prev          :   STD_ULOGIC;
 SIGNAL   DLYGL0_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL1_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL2_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL3_ipd        :   STD_ULOGIC;
 SIGNAL   DLYGL4_ipd        :   STD_ULOGIC;

 SIGNAL   GLDELAY           :   Time := 0.470 ns; -- Additional Global B Delay

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

     VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
     VitalWireDelay (DLYGL0_ipd, DLYGL0, tipd_DLYGL0);
     VitalWireDelay (DLYGL1_ipd, DLYGL1, tipd_DLYGL1);
     VitalWireDelay (DLYGL2_ipd, DLYGL2, tipd_DLYGL2);
     VitalWireDelay (DLYGL3_ipd, DLYGL3, tipd_DLYGL3);
     VitalWireDelay (DLYGL4_ipd, DLYGL4, tipd_DLYGL4);

   end block WireDelay;


  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  --
  --  get the GL output value
  --

  getGL : process(CLK_ipd, GLDELAY)

  begin

     if ( tpd_CLK_GL = VitalZeroDelay01 ) then
       GL <= transport CLK_ipd after GLDELAY;
     else
       GL <= transport CLK_ipd after VitalCalcDelay ( CLK_ipd, CLK_prev, tpd_CLK_GL );
     end if;

     CLK_prev <= CLK_ipd;

   end process getGL;

end VITAL_ACT;

configuration CFG_CLKDLYIO_VITAL of CLKDLYIO is
   for VITAL_ACT
   end for;
end CFG_CLKDLYIO_VITAL;


---- CELL PLLINT ----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
 entity PLLINT is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tpd_A_Y         : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_A          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                A               : in    STD_ULOGIC;
                Y               : out    STD_ULOGIC);
attribute VITAL_LEVEL0 of PLLINT :  entity is TRUE;
end PLLINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of PLLINT is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (A_ipd, A, tipd_A);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (A_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC is Results(1);

        -- output glitch detection variables
        VARIABLE Y_GlitchData  : VitalGlitchDataType;

        begin

           -------------------------
           --  Functionality Section
           -------------------------
        Y_zd :=TO_X01(A_ipd);


           ----------------------
           --  Path Delay Section
           ----------------------

     VitalPathDelay01 (
           OutSignal => Y,
           GlitchData => Y_GlitchData,
           OutSignalName => "Y",
           OutTemp => Y_zd,
           Paths => (
                     0 => (A_ipd'last_event,tpd_A_Y, true)),
          Mode => OnDetect,
          Xon => Xon,
          MsgOn => MsgOn,
          MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

configuration CFG_PLLINT_VITAL of PLLINT is
    for VITAL_ACT
    end for;
end CFG_PLLINT_VITAL;

---- CELL ULSICC ----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
entity ULSICC is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tipd_LSICC          : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                LSICC           : in    STD_ULOGIC);
attribute VITAL_LEVEL0 of ULSICC :  entity is TRUE;
end ULSICC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of ULSICC is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL LSICC_ipd  : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (LSICC_ipd, LSICC, tipd_LSICC);
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (LSICC_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC is Results(1);

        begin

           -------------------------
           --  Functionality Section
           -------------------------
        Y_zd :=TO_X01(LSICC_ipd);


end process;

end VITAL_ACT;

configuration CFG_ULSICC_VITAL of ULSICC is
    for VITAL_ACT
    end for;
end CFG_ULSICC_VITAL;


---- CELL ULSICC_INT ----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
entity ULSICC_INT is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tipd_USTDBY          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_LPENA           : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                USTDBY           : in    STD_ULOGIC;
                LPENA            : in    STD_ULOGIC);

attribute VITAL_LEVEL0 of ULSICC_INT :  entity is TRUE;
end ULSICC_INT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of ULSICC_INT is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL USTDBY_ipd  : STD_ULOGIC := 'X';
        SIGNAL LPENA_ipd   : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (USTDBY_ipd, USTDBY, tipd_USTDBY);
        VitalWireDelay (LPENA_ipd,  LPENA,  tipd_LPENA );
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (USTDBY_ipd, LPENA_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 downto 0)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC_VECTOR(1 downto 0) is Results(1 downto 0);

        begin

           -------------------------
           --  Functionality Section
           -------------------------
        Y_zd(0) := TO_X01(USTDBY_ipd);
        Y_zd(1) := TO_X01(LPENA_ipd);


end process;

end VITAL_ACT;

configuration CFG_ULSICC_INT_VITAL of ULSICC_INT is
    for VITAL_ACT
    end for;
end CFG_ULSICC_INT_VITAL;


---- CELL ULSICC_AUTH ----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

---- entity declaration ----
entity ULSICC_AUTH is
    generic(
                TimingChecksOn:Boolean := True;
                Xon: Boolean := False;
                InstancePath: STRING :="*";
                MsgOn: Boolean := True;
                tipd_AUTHEN          : VitalDelayType01 := (0.000 ns, 0.000 ns);
                tipd_LSICC           : VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
                AUTHEN           : in    STD_ULOGIC;
                LSICC            : in    STD_ULOGIC);

attribute VITAL_LEVEL0 of ULSICC_AUTH :  entity is TRUE;
end ULSICC_AUTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;

architecture VITAL_ACT of ULSICC_AUTH is
        attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

        SIGNAL AUTHEN_ipd  : STD_ULOGIC := 'X';
        SIGNAL LSICC_ipd   : STD_ULOGIC := 'X';

begin

        ---------------------
        --  INPUT PATH DELAYs
        ---------------------
        WireDelay : block
        begin
        VitalWireDelay (AUTHEN_ipd, AUTHEN, tipd_AUTHEN);
        VitalWireDelay (LSICC_ipd,  LSICC,  tipd_LSICC );
        end block;

        --------------------
        --  BEHAVIOR SECTION
        --------------------
        VITALBehavior : process (AUTHEN_ipd, LSICC_ipd)


        -- functionality results
        VARIABLE Results : STD_LOGIC_VECTOR(1 downto 0)  := (others => 'X');
        ALIAS Y_zd : STD_LOGIC_VECTOR(1 downto 0) is Results(1 downto 0);

        begin

           -------------------------
           --  Functionality Section
           -------------------------
        Y_zd(0) := TO_X01(AUTHEN_ipd);
        Y_zd(1) := TO_X01(LSICC_ipd);


end process;

end VITAL_ACT;

configuration CFG_ULSICC_AUTH_VITAL of ULSICC_AUTH is
    for VITAL_ACT
    end for;
end CFG_ULSICC_AUTH_VITAL;


---- CELL PLLPRIM ----
-- Timing is for the 1.5 Volt PLL - must be overwritten for the 1.2 Volt.

library IEEE;
use IEEE.std_logic_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity PLLPRIM is
  generic (
    VCOFREQUENCY       :  Real    := 0.0;
    f_CLKA_LOCK        :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

    TimingChecksOn     :  Boolean          := True;
    InstancePath       :  String           := "*";
    Xon                :  Boolean          := False;
    MsgOn              :  Boolean          := True;
    EMULATED_SYSTEM_DELAY : Time           := 3.500 ns; -- Delay Tap Additional CLK delay
    IN_DIV_DELAY          : Time           := 0.550 ns; -- Input Divider intrinsic delay
    OUT_DIV_DELAY         : Time           := 0.960 ns; -- Output Divider intrinsic delay
    MUX_DELAY             : Time           := 1.100 ns; -- MUXA/MUXB/MUXC intrinsic delay
    IN_DELAY_BYP1         : Time           := 1.523 ns; -- Input delay for CLKDIVDLY bypass mode - TIMING NOT UPDATED
    BYP_MUX_DELAY         : Time           := 0.200 ns; -- Bypass MUX intrinsic delay, not used for Ys
    GL_DRVR_DELAY         : Time           := 0.350 ns; -- Global Driver intrinsic delay
    Y_DRVR_DELAY          : Time           := 0.000 ns; -- Y Driver intrinsic delay
    FB_MUX_DELAY          : Time           := 0.900 ns; -- FBSEL MUX intrinsic delay
    X_MUX_DELAY           : Time           := 0.110 ns; -- XDLYSEL MUX intrinsic delay
    FIN_LOCK_DELAY        : Time           := 1.025 ns; -- FIN to LOCK propagation delay
    LOCK_OUT_DELAY        : Time           := 0.410 ns; -- LOCK to OUT propagation delay
    PROG_INIT_DELAY       : Time           := 1.250 ns;
    PROG_STEP_INCREMENT   : Time           := 0.360 ns;
    BYP0_CLK_GL           : Time           := 0.920 ns; -- Intrinsic delay for CLKDLY bypass mode
    CLKA_TO_REF_DELAY     : Time           := 0.600 ns;
    
    tipd_DYNSYNC       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_CLKA          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_EXTFB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_POWERDOWN     :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_CLKB          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_CLKC          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIVRST      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIVHALF     :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIVRST      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIVHALF     :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIVRST      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIVHALF     :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV5       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV6       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV5        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV6        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY2        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY3        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY4        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBSEL0        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBSEL1        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_XDLYSEL       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

    tpd_CLKA_GLA       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLA  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_GLB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_GLC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_YB        :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_YB   :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_YC        :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_YC   :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_LOCK      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_LOCK :  VitalDelayType01 := ( 0.100 ns, 0.100 ns )
   );

  port (
    DYNSYNC      : in    std_ulogic;
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    POWERDOWN    : in    std_ulogic;
    CLKB         : in    std_ulogic;
    CLKC         : in    std_ulogic;
    OADIVRST     : in    std_ulogic;
    OADIVHALF    : in    std_ulogic;
    OADIV0       : in    std_ulogic;
    OADIV1       : in    std_ulogic;
    OADIV2       : in    std_ulogic;
    OADIV3       : in    std_ulogic;
    OADIV4       : in    std_ulogic;
    OAMUX0       : in    std_ulogic;
    OAMUX1       : in    std_ulogic;
    OAMUX2       : in    std_ulogic;
    DLYGLA0      : in    std_ulogic;
    DLYGLA1      : in    std_ulogic;
    DLYGLA2      : in    std_ulogic;
    DLYGLA3      : in    std_ulogic;
    DLYGLA4      : in    std_ulogic;
    OBDIVRST     : in    std_ulogic;
    OBDIVHALF    : in    std_ulogic;
    OBDIV0       : in    std_ulogic;
    OBDIV1       : in    std_ulogic;
    OBDIV2       : in    std_ulogic;
    OBDIV3       : in    std_ulogic;
    OBDIV4       : in    std_ulogic;
    OBMUX0       : in    std_ulogic;
    OBMUX1       : in    std_ulogic;
    OBMUX2       : in    std_ulogic;
    DLYYB0       : in    std_ulogic;
    DLYYB1       : in    std_ulogic;
    DLYYB2       : in    std_ulogic;
    DLYYB3       : in    std_ulogic;
    DLYYB4       : in    std_ulogic;
    DLYGLB0      : in    std_ulogic;
    DLYGLB1      : in    std_ulogic;
    DLYGLB2      : in    std_ulogic;
    DLYGLB3      : in    std_ulogic;
    DLYGLB4      : in    std_ulogic;
    OCDIVRST     : in    std_ulogic;
    OCDIVHALF    : in    std_ulogic;
    OCDIV0       : in    std_ulogic;
    OCDIV1       : in    std_ulogic;
    OCDIV2       : in    std_ulogic;
    OCDIV3       : in    std_ulogic;
    OCDIV4       : in    std_ulogic;
    OCMUX0       : in    std_ulogic;
    OCMUX1       : in    std_ulogic;
    OCMUX2       : in    std_ulogic;
    DLYYC0       : in    std_ulogic;
    DLYYC1       : in    std_ulogic;
    DLYYC2       : in    std_ulogic;
    DLYYC3       : in    std_ulogic;
    DLYYC4       : in    std_ulogic;
    DLYGLC0      : in    std_ulogic;
    DLYGLC1      : in    std_ulogic;
    DLYGLC2      : in    std_ulogic;
    DLYGLC3      : in    std_ulogic;
    DLYGLC4      : in    std_ulogic;
    FINDIV0      : in    std_ulogic;
    FINDIV1      : in    std_ulogic;
    FINDIV2      : in    std_ulogic;
    FINDIV3      : in    std_ulogic;
    FINDIV4      : in    std_ulogic;
    FINDIV5      : in    std_ulogic;
    FINDIV6      : in    std_ulogic;
    FBDIV0       : in    std_ulogic;
    FBDIV1       : in    std_ulogic;
    FBDIV2       : in    std_ulogic;
    FBDIV3       : in    std_ulogic;
    FBDIV4       : in    std_ulogic;
    FBDIV5       : in    std_ulogic;
    FBDIV6       : in    std_ulogic;
    FBDLY0       : in    std_ulogic;
    FBDLY1       : in    std_ulogic;
    FBDLY2       : in    std_ulogic;
    FBDLY3       : in    std_ulogic;
    FBDLY4       : in    std_ulogic;
    FBSEL0       : in    std_ulogic;
    FBSEL1       : in    std_ulogic;
    XDLYSEL      : in    std_ulogic;
    VCOSEL0      : in    std_ulogic;
    VCOSEL1      : in    std_ulogic;
    VCOSEL2      : in    std_ulogic;
    GLA          : out   std_ulogic;
    LOCK         : out   std_ulogic;
    GLB          : out   std_ulogic;
    YB           : out   std_ulogic;
    GLC          : out   std_ulogic;
    YC           : out   std_ulogic
   );

  attribute VITAL_LEVEL0 of PLLPRIM : entity is TRUE;
end PLLPRIM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of PLLPRIM is
attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal DYNSYNC_ipd            : std_ulogic;
  signal CLKA_ipd               : std_ulogic;
  signal EXTFB_ipd              : std_ulogic;
  signal POWERDOWN_ipd          : std_ulogic;
  signal CLKB_ipd               : std_ulogic;
  signal CLKC_ipd               : std_ulogic;
  signal OADIVRST_ipd           : std_ulogic;
  signal OADIVHALF_ipd          : std_ulogic;
  signal OADIV0_ipd             : std_ulogic;
  signal OADIV1_ipd             : std_ulogic;
  signal OADIV2_ipd             : std_ulogic;
  signal OADIV3_ipd             : std_ulogic;
  signal OADIV4_ipd             : std_ulogic;
  signal OAMUX0_ipd             : std_ulogic;
  signal OAMUX1_ipd             : std_ulogic;
  signal OAMUX2_ipd             : std_ulogic;
  signal DLYGLA0_ipd            : std_ulogic;
  signal DLYGLA1_ipd            : std_ulogic;
  signal DLYGLA2_ipd            : std_ulogic;
  signal DLYGLA3_ipd            : std_ulogic;
  signal DLYGLA4_ipd            : std_ulogic;
  signal OBDIVRST_ipd           : std_ulogic;
  signal OBDIVHALF_ipd          : std_ulogic;
  signal OBDIV0_ipd             : std_ulogic;
  signal OBDIV1_ipd             : std_ulogic;
  signal OBDIV2_ipd             : std_ulogic;
  signal OBDIV3_ipd             : std_ulogic;
  signal OBDIV4_ipd             : std_ulogic;
  signal OBMUX0_ipd             : std_ulogic;
  signal OBMUX1_ipd             : std_ulogic;
  signal OBMUX2_ipd             : std_ulogic;
  signal DLYYB0_ipd             : std_ulogic;
  signal DLYYB1_ipd             : std_ulogic;
  signal DLYYB2_ipd             : std_ulogic;
  signal DLYYB3_ipd             : std_ulogic;
  signal DLYYB4_ipd             : std_ulogic;
  signal DLYGLB0_ipd            : std_ulogic;
  signal DLYGLB1_ipd            : std_ulogic;
  signal DLYGLB2_ipd            : std_ulogic;
  signal DLYGLB3_ipd            : std_ulogic;
  signal DLYGLB4_ipd            : std_ulogic;
  signal OCDIVRST_ipd           : std_ulogic;
  signal OCDIVHALF_ipd          : std_ulogic;
  signal OCDIV0_ipd             : std_ulogic;
  signal OCDIV1_ipd             : std_ulogic;
  signal OCDIV2_ipd             : std_ulogic;
  signal OCDIV3_ipd             : std_ulogic;
  signal OCDIV4_ipd             : std_ulogic;
  signal OCMUX0_ipd             : std_ulogic;
  signal OCMUX1_ipd             : std_ulogic;
  signal OCMUX2_ipd             : std_ulogic;
  signal DLYYC0_ipd             : std_ulogic;
  signal DLYYC1_ipd             : std_ulogic;
  signal DLYYC2_ipd             : std_ulogic;
  signal DLYYC3_ipd             : std_ulogic;
  signal DLYYC4_ipd             : std_ulogic;
  signal DLYGLC0_ipd            : std_ulogic;
  signal DLYGLC1_ipd            : std_ulogic;
  signal DLYGLC2_ipd            : std_ulogic;
  signal DLYGLC3_ipd            : std_ulogic;
  signal DLYGLC4_ipd            : std_ulogic;
  signal FINDIV0_ipd            : std_ulogic;
  signal FINDIV1_ipd            : std_ulogic;
  signal FINDIV2_ipd            : std_ulogic;
  signal FINDIV3_ipd            : std_ulogic;
  signal FINDIV4_ipd            : std_ulogic;
  signal FINDIV5_ipd            : std_ulogic;
  signal FINDIV6_ipd            : std_ulogic;
  signal FBDIV0_ipd             : std_ulogic;
  signal FBDIV1_ipd             : std_ulogic;
  signal FBDIV2_ipd             : std_ulogic;
  signal FBDIV3_ipd             : std_ulogic;
  signal FBDIV4_ipd             : std_ulogic;
  signal FBDIV5_ipd             : std_ulogic;
  signal FBDIV6_ipd             : std_ulogic;
  signal FBDLY0_ipd             : std_ulogic;
  signal FBDLY1_ipd             : std_ulogic;
  signal FBDLY2_ipd             : std_ulogic;
  signal FBDLY3_ipd             : std_ulogic;
  signal FBDLY4_ipd             : std_ulogic;
  signal FBSEL0_ipd             : std_ulogic;
  signal FBSEL1_ipd             : std_ulogic;
  signal XDLYSEL_ipd            : std_ulogic;
  signal VCOSEL0_ipd            : std_ulogic;
  signal VCOSEL1_ipd            : std_ulogic;
  signal VCOSEL2_ipd            : std_ulogic;

  signal AOUT                   : std_logic := 'X';
  signal BOUT                   : std_logic := 'X';
  signal COUT                   : std_logic := 'X';

  signal PLLCLK                 : std_logic := 'X';      -- PLL Core Output Clock 
                                                         -- with DIVN and DIVM applied
  signal CLKA_period            : Time      := 0.000 ns; -- Current CLKA period

  signal PLLCLK_pw              : Time      := 10.0 ns; -- PLLCLK pulse width
  signal PLLCLK_period          : Time      := 10.0 ns;

  signal DIVN                   : Integer := 1; -- Divide by N divisor - range 1 to 128
  signal DIVM                   : Integer := 1; -- Multiply by M multiplier - range 1 to 128
  signal DIVU                   : Integer := 1; -- Divide by U divisor - range 1 to 32
  signal DIVV                   : Integer := 1; -- Divide by V divisor - range 1 to 32
  signal DIVW                   : Integer := 1; -- Divide by W divisor - range 1 to 32
  signal fb_loop_div            : Integer := 1; -- Total division of feedback loop

  signal halveA                 : std_logic := 'X';
  signal halveB                 : std_logic := 'X';
  signal halveC                 : std_logic := 'X';

  signal CLKA2X                 : std_logic := 'X';
  signal CLKB2X                 : std_logic := 'X';
  signal CLKC2X                 : std_logic := 'X';

  signal UIN                    : std_logic := 'X'; -- Output of MUXA
  signal VIN                    : std_logic := 'X'; -- Output of MUXB
  signal WIN                    : std_logic := 'X'; -- Output of MUXC

  signal FBDELAY                : Time := 0.000 ns; -- Feedback delay
  signal DTDELAY                : Time := 0.000 ns; -- Delay Tap delay
  signal PLLDELAY               : Time := 0.000 ns; -- Sum of Feedback and Delay Tap delays
  signal YBDELAY                : Time := 0.000 ns; -- Additional Global B Delay
  signal GLBDELAY               : Time := 0.000 ns; -- Additional Global B Delay
  signal YCDELAY                : Time := 0.000 ns; -- Additional Global C Delay
  signal GLCDELAY               : Time := 0.000 ns; -- Additional Global C Delay
  signal GLADELAY               : Time := 0.000 ns; -- Additional Global A Delay

  signal FBSEL                  : std_logic_vector( 1 downto 0 ) := "XX";
  signal FBSEL_illegal          : Boolean := False; -- True when FBSEL = 00

  signal OAMUX_config           : integer := -1;
  signal OBMUX_config           : integer := -1;
  signal OCMUX_config           : integer := -1;

  signal internal_lock          : boolean   := false;
  signal fin_period             : Time      := 0.000 ns;
  signal extfbin_fin_drift      : time      := 0 ps;
  signal locked                 : std_logic := '0'; -- 1 when PLL is externally locked as well as internally locked
  signal locked_vco0_edges      : integer   := -1;
  signal vco0_divu              : std_logic := '0';
  signal vco0_divv              : std_logic := '0';
  signal vco0_divw              : std_logic := '0';
  signal fin                    : std_logic := '0';
  signal CLKA_period_stable     : boolean   := false;

  signal using_EXTFB            : std_logic := 'X';
  signal EXTFB_delay_dtrmd      : Boolean   := false;
  signal calibrate_EXTFB_delay  : std_logic := '0';
  signal GLA_free_running       : std_logic := '1';
  signal AOUT_using_EXTFB       : std_logic := '1';
  signal GLA_pw                 : time      := 10.0 ns; -- Only used for external feedback
  signal GLA_EXTFB_rise_dly     : time      := 0.0 ns;  -- Only meaningful for external feedback
  signal GLA_EXTFB_fall_dly     : time      := 0.0 ns;  -- Only meaningful for external feedback
  signal EXTFB_period           : time      := 20.0 ns;  -- Only meaningful for external feedback
  signal expected_EXTFB         : std_logic := 'X';
  signal external_dly_correct   : std_logic := 'X';

  signal gla_muxed_delay        : time      := 0.000 ns;
  signal glb_muxed_delay        : time      := 0.000 ns;
  signal glc_muxed_delay        : time      := 0.000 ns;

  signal internal_fb_delay      : time      := 0.000 ns;
  signal external_fb_delay      : time      := 0.000 ns;
  signal normalized_fb_delay    : time      := 0.000 ns; -- Sum of all delays in the feedback loop from VCO to FBIN normalized to be less than or equal to fin period so that no negative delay assignments are made.

  signal CLKA_2_GLA_dly         : time      := 0.000 ns;
  signal CLKA_2_GLA_bypass0_dly : time      := 0.000 ns;
  signal CLKA_2_GLA_bypass1_dly : time      := 0.000 ns;
  signal CLKA_2_GLB_dly         : time      := 0.000 ns;
  signal CLKB_2_GLB_bypass0_dly : time      := 0.000 ns;
  signal CLKB_2_GLB_bypass1_dly : time      := 0.000 ns;
  signal CLKA_2_YB_dly          : time      := 0.000 ns;
  signal CLKB_2_YB_bypass1_dly  : time      := 0.000 ns;
  signal CLKA_2_GLC_dly         : time      := 0.000 ns;
  signal CLKC_2_GLC_bypass0_dly : time      := 0.000 ns;
  signal CLKC_2_GLC_bypass1_dly : time      := 0.000 ns;
  signal CLKA_2_YC_dly          : time      := 0.000 ns;
  signal CLKC_2_YC_bypass1_dly  : time      := 0.000 ns;
  signal CLKA_2_LOCK_dly        : time      := 0.000 ns;


  -- Use this instead of CONV_INTEGER to avoid ambiguous warnings
  function ulogic2int(
    vec  : std_ulogic_vector )
    return integer is
    variable result : integer;
    variable i : integer;
  begin
    result := 0;
    for i in vec'range loop
      result := result * 2;
      if vec(i) = '1' then
        result := result + 1;
      end if;
    end loop;
    return result;
  end function ulogic2int;

  function output_mux_delay( 
    outmux      : integer;
    vcobit2     : std_logic;
    vcobit1     : std_logic;
    fbdly_delay : time;
    vco_pw      : time )
    return time is
    variable result : time;
  begin
     case outmux is
        when 1  => result := IN_DELAY_BYP1;
        when 2  => result := MUX_DELAY + fbdly_delay;
        when 5  => if ( ( vcobit2 = '1') and ( vcobit1 = '1') ) then
                         result := MUX_DELAY + ( vco_pw / 2.0 );
                       else
                         result := MUX_DELAY + ( vco_pw * 1.5 );
                       end if;
        when 6  => result := MUX_DELAY + vco_pw;
        when 7  => if ( ( vcobit2 = '1') and ( vcobit1 = '1') ) then
                         result := MUX_DELAY + ( vco_pw * 1.5 );
                       else
                         result := MUX_DELAY + ( vco_pw / 2.0 );
                       end if;
        when others => result := MUX_DELAY;
     end case;
     return result;
  end function output_mux_delay;


  function output_mux_driver( 
    outmux      : integer;
    halved      : std_logic;
    bypass      : std_logic;
    bypass2x    : std_logic;
    vco         : std_logic )
    return std_logic is
    variable result : std_logic;
  begin
     case outmux is
        when 1  => if ( '1' = halved ) then
                          result := bypass2x;
                       elsif ( '0' = halved ) then
                          result := bypass;
                       else
                          result := 'X';
                       end if;
        when 2  => result := vco;
        when 4  => result := vco;
        when 5  => result := vco;
        when 6  => result := vco;
        when 7  => result := vco;
        when others => result := 'X';
     end case;
     return result;
  end function output_mux_driver;

  begin

    ---------------------
    --  INPUT PATH DELAYs
    ---------------------
    WireDelay : block

    begin

      VitalWireDelay ( DYNSYNC_ipd,   DYNSYNC,   tipd_DYNSYNC   );
      VitalWireDelay ( CLKA_ipd,      CLKA,      tipd_CLKA      );
      VitalWireDelay ( EXTFB_ipd,     EXTFB,     tipd_EXTFB     );
      VitalWireDelay ( POWERDOWN_ipd, POWERDOWN, tipd_POWERDOWN );
      VitalWireDelay ( CLKB_ipd,      CLKB,      tipd_CLKB      );
      VitalWireDelay ( CLKC_ipd,      CLKC,      tipd_CLKC      );
      VitalWireDelay ( OADIVRST_ipd,  OADIVRST,  tipd_OADIVRST  );
      VitalWireDelay ( OADIVHALF_ipd, OADIVHALF, tipd_OADIVHALF );
      VitalWireDelay ( OADIV0_ipd,    OADIV0,    tipd_OADIV0    );
      VitalWireDelay ( OADIV1_ipd,    OADIV1,    tipd_OADIV1    );
      VitalWireDelay ( OADIV2_ipd,    OADIV2,    tipd_OADIV2    );
      VitalWireDelay ( OADIV3_ipd,    OADIV3,    tipd_OADIV3    );
      VitalWireDelay ( OADIV4_ipd,    OADIV4,    tipd_OADIV4    );
      VitalWireDelay ( OAMUX0_ipd,    OAMUX0,    tipd_OAMUX0    );
      VitalWireDelay ( OAMUX1_ipd,    OAMUX1,    tipd_OAMUX1    );
      VitalWireDelay ( OAMUX2_ipd,    OAMUX2,    tipd_OAMUX2    );
      VitalWireDelay ( DLYGLA0_ipd,   DLYGLA0,   tipd_DLYGLA0   );
      VitalWireDelay ( DLYGLA1_ipd,   DLYGLA1,   tipd_DLYGLA1   );
      VitalWireDelay ( DLYGLA2_ipd,   DLYGLA2,   tipd_DLYGLA2   );
      VitalWireDelay ( DLYGLA3_ipd,   DLYGLA3,   tipd_DLYGLA3   );
      VitalWireDelay ( DLYGLA4_ipd,   DLYGLA4,   tipd_DLYGLA4   );
      VitalWireDelay ( OBDIVRST_ipd,  OBDIVRST,  tipd_OBDIVRST  );
      VitalWireDelay ( OBDIVHALF_ipd, OBDIVHALF, tipd_OBDIVHALF );
      VitalWireDelay ( OBDIV0_ipd,    OBDIV0,    tipd_OBDIV0    );
      VitalWireDelay ( OBDIV1_ipd,    OBDIV1,    tipd_OBDIV1    );
      VitalWireDelay ( OBDIV2_ipd,    OBDIV2,    tipd_OBDIV2    );
      VitalWireDelay ( OBDIV3_ipd,    OBDIV3,    tipd_OBDIV3    );
      VitalWireDelay ( OBDIV4_ipd,    OBDIV4,    tipd_OBDIV4    );
      VitalWireDelay ( OBMUX0_ipd,    OBMUX0,    tipd_OBMUX0    );
      VitalWireDelay ( OBMUX1_ipd,    OBMUX1,    tipd_OBMUX1    );
      VitalWireDelay ( OBMUX2_ipd,    OBMUX2,    tipd_OBMUX2    );
      VitalWireDelay ( DLYYB0_ipd,    DLYYB0,    tipd_DLYYB0    );
      VitalWireDelay ( DLYYB1_ipd,    DLYYB1,    tipd_DLYYB1    );
      VitalWireDelay ( DLYYB2_ipd,    DLYYB2,    tipd_DLYYB2    );
      VitalWireDelay ( DLYYB3_ipd,    DLYYB3,    tipd_DLYYB3    );
      VitalWireDelay ( DLYYB4_ipd,    DLYYB4,    tipd_DLYYB4    );
      VitalWireDelay ( DLYGLB0_ipd,   DLYGLB0,   tipd_DLYGLB0   );
      VitalWireDelay ( DLYGLB1_ipd,   DLYGLB1,   tipd_DLYGLB1   );
      VitalWireDelay ( DLYGLB2_ipd,   DLYGLB2,   tipd_DLYGLB2   );
      VitalWireDelay ( DLYGLB3_ipd,   DLYGLB3,   tipd_DLYGLB3   );
      VitalWireDelay ( DLYGLB4_ipd,   DLYGLB4,   tipd_DLYGLB4   );
      VitalWireDelay ( OCDIVRST_ipd,  OCDIVRST,  tipd_OCDIVRST  );
      VitalWireDelay ( OCDIVHALF_ipd, OCDIVHALF, tipd_OCDIVHALF );
      VitalWireDelay ( OCDIV0_ipd,    OCDIV0,    tipd_OCDIV0    );
      VitalWireDelay ( OCDIV1_ipd,    OCDIV1,    tipd_OCDIV1    );
      VitalWireDelay ( OCDIV2_ipd,    OCDIV2,    tipd_OCDIV2    );
      VitalWireDelay ( OCDIV3_ipd,    OCDIV3,    tipd_OCDIV3    );
      VitalWireDelay ( OCDIV4_ipd,    OCDIV4,    tipd_OCDIV4    );
      VitalWireDelay ( OCMUX0_ipd,    OCMUX0,    tipd_OCMUX0    );
      VitalWireDelay ( OCMUX1_ipd,    OCMUX1,    tipd_OCMUX1    );
      VitalWireDelay ( OCMUX2_ipd,    OCMUX2,    tipd_OCMUX2    );
      VitalWireDelay ( DLYYC0_ipd,    DLYYC0,    tipd_DLYYC0    );
      VitalWireDelay ( DLYYC1_ipd,    DLYYC1,    tipd_DLYYC1    );
      VitalWireDelay ( DLYYC2_ipd,    DLYYC2,    tipd_DLYYC2    );
      VitalWireDelay ( DLYYC3_ipd,    DLYYC3,    tipd_DLYYC3    );
      VitalWireDelay ( DLYYC4_ipd,    DLYYC4,    tipd_DLYYC4    );
      VitalWireDelay ( DLYGLC0_ipd,   DLYGLC0,   tipd_DLYGLC0   );
      VitalWireDelay ( DLYGLC1_ipd,   DLYGLC1,   tipd_DLYGLC1   );
      VitalWireDelay ( DLYGLC2_ipd,   DLYGLC2,   tipd_DLYGLC2   );
      VitalWireDelay ( DLYGLC3_ipd,   DLYGLC3,   tipd_DLYGLC3   );
      VitalWireDelay ( DLYGLC4_ipd,   DLYGLC4,   tipd_DLYGLC4   );
      VitalWireDelay ( FINDIV0_ipd,   FINDIV0,   tipd_FINDIV0   );
      VitalWireDelay ( FINDIV1_ipd,   FINDIV1,   tipd_FINDIV1   );
      VitalWireDelay ( FINDIV2_ipd,   FINDIV2,   tipd_FINDIV2   );
      VitalWireDelay ( FINDIV3_ipd,   FINDIV3,   tipd_FINDIV3   );
      VitalWireDelay ( FINDIV4_ipd,   FINDIV4,   tipd_FINDIV4   );
      VitalWireDelay ( FINDIV5_ipd,   FINDIV5,   tipd_FINDIV5   );
      VitalWireDelay ( FINDIV6_ipd,   FINDIV6,   tipd_FINDIV6   );
      VitalWireDelay ( FBDIV0_ipd,    FBDIV0,    tipd_FBDIV0    );
      VitalWireDelay ( FBDIV1_ipd,    FBDIV1,    tipd_FBDIV1    );
      VitalWireDelay ( FBDIV2_ipd,    FBDIV2,    tipd_FBDIV2    );
      VitalWireDelay ( FBDIV3_ipd,    FBDIV3,    tipd_FBDIV3    );
      VitalWireDelay ( FBDIV4_ipd,    FBDIV4,    tipd_FBDIV4    );
      VitalWireDelay ( FBDIV5_ipd,    FBDIV5,    tipd_FBDIV5    );
      VitalWireDelay ( FBDIV6_ipd,    FBDIV6,    tipd_FBDIV6    );
      VitalWireDelay ( FBDLY0_ipd,    FBDLY0,    tipd_FBDLY0    );
      VitalWireDelay ( FBDLY1_ipd,    FBDLY1,    tipd_FBDLY1    );
      VitalWireDelay ( FBDLY2_ipd,    FBDLY2,    tipd_FBDLY2    );
      VitalWireDelay ( FBDLY3_ipd,    FBDLY3,    tipd_FBDLY3    );
      VitalWireDelay ( FBDLY4_ipd,    FBDLY4,    tipd_FBDLY4    );
      VitalWireDelay ( FBSEL0_ipd,    FBSEL0,    tipd_FBSEL0    );
      VitalWireDelay ( FBSEL1_ipd,    FBSEL1,    tipd_FBSEL1    );
      VitalWireDelay ( XDLYSEL_ipd,   XDLYSEL,   tipd_XDLYSEL   );
      VitalWireDelay ( VCOSEL0_ipd,   VCOSEL0,   tipd_VCOSEL0   );
      VitalWireDelay ( VCOSEL1_ipd,   VCOSEL1,   tipd_VCOSEL1   );
      VitalWireDelay ( VCOSEL2_ipd,   VCOSEL2,   tipd_VCOSEL2   );
 
    end block WireDelay;

    -- #########################################################
    -- # Behavior Section
    -- #########################################################

    OAMUX_config <= ulogic2int( OAMUX2_ipd & OAMUX1_ipd & OAMUX0_ipd );
    OBMUX_config <= ulogic2int( OBMUX2_ipd & OBMUX1_ipd & OBMUX0_ipd );
    OCMUX_config <= ulogic2int( OCMUX2_ipd & OCMUX1_ipd & OCMUX0_ipd );
    FBSEL <= TO_X01( FBSEL1_ipd & FBSEL0_ipd );

    CLKA_2_GLA_dly         <= CLKA_TO_REF_DELAY + IN_DIV_DELAY + fin_period - normalized_fb_delay + gla_muxed_delay + OUT_DIV_DELAY + BYP_MUX_DELAY + GLADELAY + GL_DRVR_DELAY;
    CLKA_2_GLA_bypass0_dly <= BYP0_CLK_GL + GLADELAY;
    CLKA_2_GLA_bypass1_dly <= gla_muxed_delay + OUT_DIV_DELAY + BYP_MUX_DELAY + GLADELAY + GL_DRVR_DELAY;

    CLKA_2_GLB_dly         <= CLKA_TO_REF_DELAY + IN_DIV_DELAY + fin_period - normalized_fb_delay + glb_muxed_delay + OUT_DIV_DELAY + BYP_MUX_DELAY + GLBDELAY + GL_DRVR_DELAY;
    CLKB_2_GLB_bypass0_dly <= BYP0_CLK_GL + GLBDELAY;
    CLKB_2_GLB_bypass1_dly <= glb_muxed_delay + OUT_DIV_DELAY + BYP_MUX_DELAY + GLBDELAY + GL_DRVR_DELAY;
    CLKA_2_YB_dly          <= CLKA_TO_REF_DELAY + IN_DIV_DELAY + fin_period - normalized_fb_delay + glb_muxed_delay + OUT_DIV_DELAY + YBDELAY + Y_DRVR_DELAY;
    CLKB_2_YB_bypass1_dly  <= glb_muxed_delay + OUT_DIV_DELAY + YBDELAY + Y_DRVR_DELAY;

    CLKA_2_GLC_dly         <= CLKA_TO_REF_DELAY + IN_DIV_DELAY + fin_period - normalized_fb_delay + glc_muxed_delay + OUT_DIV_DELAY + BYP_MUX_DELAY + GLCDELAY + GL_DRVR_DELAY;
    CLKC_2_GLC_bypass0_dly <= BYP0_CLK_GL + GLCDELAY;
    CLKC_2_GLC_bypass1_dly <= glc_muxed_delay + OUT_DIV_DELAY + BYP_MUX_DELAY + GLCDELAY + GL_DRVR_DELAY;
    CLKA_2_YC_dly          <= CLKA_TO_REF_DELAY + IN_DIV_DELAY + fin_period - normalized_fb_delay + glc_muxed_delay + OUT_DIV_DELAY + YCDELAY + Y_DRVR_DELAY;
    CLKC_2_YC_bypass1_dly  <= glc_muxed_delay + OUT_DIV_DELAY + YCDELAY + Y_DRVR_DELAY;

    CLKA_2_LOCK_dly        <= CLKA_TO_REF_DELAY + IN_DIV_DELAY + fin_period - normalized_fb_delay + LOCK_OUT_DELAY;

    delay_LOCK: process( locked )
    begin
       if ( '1' = locked ) then
          LOCK <= transport locked after CLKA_2_LOCK_dly;
       else
          LOCK <= locked;
       end if;
    end process delay_LOCK;

    Deskew : process ( XDLYSEL_ipd )
      variable DelayVal             : Time := 0.000 ns;
    begin
      if (XDLYSEL_ipd = '1') then
        DelayVal := EMULATED_SYSTEM_DELAY;
      else
        DelayVal := 0.0 ns;
      end if;
      DTDELAY <= DelayVal;
    end process Deskew;

    GetFBDelay : process ( FBDLY0_ipd, FBDLY1_ipd, FBDLY2_ipd, FBDLY3_ipd, FBDLY4_ipd )
      variable step : integer;
    begin
      step := ulogic2int( FBDLY4_ipd & FBDLY3_ipd & FBDLY2_ipd & FBDLY1_ipd & FBDLY0_ipd );
      FBDELAY <= ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
    end process GetFBDelay;

    GetGLBDelay : process ( DLYGLB0_ipd, DLYGLB1_ipd, DLYGLB2_ipd, DLYGLB3_ipd, DLYGLB4_ipd )
      variable step : integer;
    begin
      step := ulogic2int( DLYGLB4_ipd & DLYGLB3_ipd & DLYGLB2_ipd & DLYGLB1_ipd & DLYGLB0_ipd );
      if ( step = 0 ) then
        GLBDELAY <= 0.0 ns;
      else
        GLBDELAY <= ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
      end if;
    end process GetGLBDelay;

    GetYBDelay : process ( DLYYB0_ipd, DLYYB1_ipd, DLYYB2_ipd, DLYYB3_ipd, DLYYB4_ipd )
      variable step : integer;
    begin
      step := ulogic2int( DLYYB4_ipd & DLYYB3_ipd & DLYYB2_ipd & DLYYB1_ipd & DLYYB0_ipd );
      YBDELAY <= ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
    end process GetYBDelay;

    GetGLCDelay : process ( DLYGLC0_ipd, DLYGLC1_ipd, DLYGLC2_ipd, DLYGLC3_ipd, DLYGLC4_ipd )
      variable step : integer;
    begin
      step := ulogic2int( DLYGLC4_ipd & DLYGLC3_ipd & DLYGLC2_ipd & DLYGLC1_ipd & DLYGLC0_ipd );
      if ( step = 0 ) then
        GLCDELAY <= 0.0 ns;
      else
        GLCDELAY <= ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
      end if;
    end process GetGLCDelay;

    GetYCDelay : process ( DLYYC0_ipd, DLYYC1_ipd, DLYYC2_ipd, DLYYC3_ipd, DLYYC4_ipd )
      variable step : integer;
    begin
      step := ulogic2int( DLYYC4_ipd & DLYYC3_ipd & DLYYC2_ipd & DLYYC1_ipd & DLYYC0_ipd );
      YCDELAY <= ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
    end process GetYCDelay;

    GetGLADelay : process ( DLYGLA0_ipd, DLYGLA1_ipd, DLYGLA2_ipd, DLYGLA3_ipd, DLYGLA4_ipd )
      variable step : integer;
    begin
      step := ulogic2int( DLYGLA4_ipd & DLYGLA3_ipd & DLYGLA2_ipd & DLYGLA1_ipd & DLYGLA0_ipd );
      if ( step = 0 ) then
        GLADELAY <= 0.0 ns;
      else
        GLADELAY <= ( step * PROG_STEP_INCREMENT ) + PROG_INIT_DELAY;
      end if;
    end process GetGLADelay;

    DIVM <= ulogic2int( FBDIV6_ipd & FBDIV5_ipd & FBDIV4_ipd & FBDIV3_ipd & 
                        FBDIV2_ipd & FBDIV1_ipd & FBDIV0_ipd ) + 1;

    DIVN <= ulogic2int( FINDIV6_ipd & FINDIV5_ipd & FINDIV4_ipd & FINDIV3_ipd & 
                        FINDIV2_ipd & FINDIV1_ipd & FINDIV0_ipd ) + 1;

    DIVU <= ulogic2int( OADIV4_ipd & OADIV3_ipd & OADIV2_ipd & OADIV1_ipd & OADIV0_ipd ) + 1;

    DIVV <= ulogic2int( OBDIV4_ipd & OBDIV3_ipd & OBDIV2_ipd & OBDIV1_ipd & OBDIV0_ipd ) + 1;

    DIVW <= ulogic2int( OCDIV4_ipd & OCDIV3_ipd & OCDIV2_ipd & OCDIV1_ipd & OCDIV0_ipd ) + 1;

    check_OADIVHALF : process
    begin
       wait on OADIVHALF_ipd, DIVU, OAMUX_config;
       if ( '1' = TO_X01( OADIVHALF_ipd ) ) then
         if ( 1 /= OAMUX_config ) then
            assert false
               report "Illegal configuration.  OADIVHALF can only be used when OAMUX = 001. OADIVHALF ignored."
               severity warning;
            halveA <= '0';
         elsif ( ( DIVU < 3 ) or ( DIVU > 29 ) or ( ( DIVU mod 2 ) /= 1 ) ) then
            assert false
               report "Illegal configuration. Only even OADIV values from 2 to 28 (inclusive) are allowed with OADIVHALF."
               severity warning;
            halveA <= 'X';
         else
            halveA <= '1';
         end if;
       elsif ( OADIVHALF_ipd'event and ( 'X' = TO_X01( OADIVHALF_ipd ) ) ) then
          assert false
             report "OADIVHALF unknown."
             severity warning;
          halveA <= 'X';
       else
          halveA <= '0';
       end if;
    end process check_OADIVHALF;

    check_OBDIVHALF : process
    begin
       wait on OBDIVHALF_ipd, DIVV, OBMUX_config;
       if ( '1' = TO_X01( OBDIVHALF_ipd ) ) then
         if ( 1 /= OBMUX_config ) then
            assert false
               report "Illegal configuration.  OBDIVHALF can only be used when OBMUX = 001. OBDIVHALF ignored."
               severity warning;
            halveB <= '0';
         elsif ( ( DIVV < 3 ) or ( DIVV > 29 ) or ( ( DIVV mod 2 ) /= 1 ) ) then
            assert false
               report "Illegal configuration. Only even OBDIV values from 2 to 28 (inclusive) are allowed with OBDIVHALF."
               severity warning;
            halveB <= 'X';
         else
            halveB <= '1';
         end if;
       elsif ( OBDIVHALF_ipd'event and ( 'X' = TO_X01( OBDIVHALF_ipd ) ) ) then
          assert false
             report "OBDIVHALF unknown."
             severity warning;
          halveB <= 'X';
       else
          halveB <= '0';
       end if;
    end process check_OBDIVHALF;

    check_OCDIVHALF : process
    begin
       wait on OCDIVHALF_ipd, DIVW, OCMUX_config;
       if ( '1' = TO_X01( OCDIVHALF_ipd ) ) then
         if ( 1 /= OCMUX_config ) then
            assert false
               report "Illegal configuration.  OCDIVHALF can only be used when OCMUX = 001. OCDIVHALF ignored."
               severity warning;
            halveC <= '0';
         elsif ( ( DIVW < 3 ) or ( DIVW > 29 ) or ( ( DIVW mod 2 ) /= 1 ) ) then
            assert false
               report "Illegal configuration. Only even OCDIV values from 2 to 28 (inclusive) are allowed with OCDIVHALF."
               severity warning;
            halveC <= 'X';
         else
            halveC <= '1';
         end if;
       elsif ( OCDIVHALF_ipd'event and ( 'X' = TO_X01( OCDIVHALF_ipd ) ) ) then
          assert false
             report "OCDIVHALF unknown."
             severity warning;
          halveC <= 'X';
       else
          halveC <= '0';
       end if;
    end process check_OCDIVHALF;

    gla_muxed_delay <= output_mux_delay( OAMUX_config, VCOSEL2_ipd, VCOSEL1_ipd, FBDELAY, PLLCLK_pw );
    glb_muxed_delay <= output_mux_delay( OBMUX_config, VCOSEL2_ipd, VCOSEL1_ipd, FBDELAY, PLLCLK_pw );
    glc_muxed_delay <= output_mux_delay( OCMUX_config, VCOSEL2_ipd, VCOSEL1_ipd, FBDELAY, PLLCLK_pw );

    get_internal_fb_dly : process( FBSEL, FBDELAY, DTDELAY, fin_period )
       variable fb_delay : time;
    begin
       fb_delay := IN_DIV_DELAY + X_MUX_DELAY + DTDELAY + FB_MUX_DELAY;
       if ( "10" = FBSEL ) then
         fb_delay := fb_delay + FBDELAY;
       end if;
       internal_fb_delay <= fb_delay;
    end process get_internal_fb_dly;

    external_fb_delay <= IN_DIV_DELAY + X_MUX_DELAY + DTDELAY + FB_MUX_DELAY + GL_DRVR_DELAY + GLADELAY + BYP_MUX_DELAY + OUT_DIV_DELAY + gla_muxed_delay + GLA_EXTFB_rise_dly;

    normalize_fb_dly : process( using_EXTFB, internal_fb_delay, external_fb_delay, fin_period )
       variable norm : time;
    begin
       if ( using_EXTFB = '1' ) then
          norm := external_fb_delay;
       else
          norm := internal_fb_delay;
       end if;
       if ( 0 ns >= fin_period ) then
          norm := 0 ns;
       else
         while ( norm > fin_period ) loop
            norm := norm - fin_period;
         end loop;
       end if;
       normalized_fb_delay <= norm;
    end process normalize_fb_dly;

    check_FBSEL : process
    begin
      wait on FBSEL, OAMUX_config, OBMUX_config, OCMUX_config, DIVM, DIVU, DIVN, CLKA_period_stable, PLLCLK_period, external_fb_delay;
      if ( IS_X( FBSEL ) ) then
         FBSEL_illegal <= true;
         assert ( not FBSEL'event )
            report "Warning: FBSEL is unknown." 
            severity Warning;
      elsif ( "00" = FBSEL ) then -- Grounded.
         FBSEL_illegal <= true;
         assert ( not FBSEL'event )
            report "Warning: Illegal FBSEL configuration 00." 
            severity Warning;
      elsif ( "11" = FBSEL ) then -- External feedback
         if ( 2 > OAMUX_config ) then
            FBSEL_illegal <= true;
            assert  ( not ( FBSEL'event or OAMUX_config'event ) )
               report "Illegal configuration. GLA cannot be in bypass mode (OAMUX = 000 or OAMUX = 001) when using external feedback (FBSEL = 11)." 
               severity Warning;
         elsif ( DIVM < 5 ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or DIVM'event ) )
               report "Error: FBDIV must be greater than 4 when using external feedback (FBSEL = 11)."
               severity Error;
         elsif ( ( DIVM * DIVU ) > 232 ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or DIVM'event or DIVU'event ) )
               report "Error: Product of FBDIV and OADIV must be less than 233 when using external feedback (FBSEL = 11)."
               severity Error;
         elsif ( ( DIVN mod DIVU ) /= 0 ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or DIVN'event or DIVU'event ) )
               report "Error: Division factor FINDIV must be a multiple of OADIV when using external feedback (FBSEL = 11)."
               severity Error;
         elsif ( CLKA_period_stable and EXTFB_delay_dtrmd and
                 ( ( 1 < OBMUX_config ) or ( 1 < OCMUX_config ) ) and
                 ( ( external_fb_delay >= CLKA_period ) or ( external_fb_delay >= PLLCLK_period ) ) ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or CLKA_period_stable'event or external_fb_delay'event or PLLCLK_period'event ) )
              report "Error: Total sum of delays in the feedback path must be less than 1 VCO period AND less than 1 CLKA period when V and/or W dividers when using external feedback (FBSEL = 11)."
               severity Error;
         else
            FBSEL_illegal <= false;
         end if;
      else
         FBSEL_illegal <= false;
      end if;
    end process check_FBSEL;

    -- Mimicing silicon - no need for a 50/50 duty cycle and this way fin only changes on rising edge of CLKA (except when DIVN is 1)
    gen_fin: process
      variable num_CLKA_re   : integer;
    begin
       wait until rising_edge( CLKA_ipd );
       fin <= '1';
       num_CLKA_re := 0;
       while ( 'X' /= TO_X01( CLKA_ipd ) ) loop
          wait on CLKA_ipd;
          if ( 1 = DIVN )then
             fin <= CLKA_ipd;
          elsif ( '1' = CLKA_ipd ) then
             num_CLKA_re := num_CLKA_re + 1;
             if ( ( num_CLKA_re mod DIVN  ) = 0 ) then
                fin <= '1';
                num_CLKA_re := 0;
             elsif ( ( num_CLKA_re mod DIVN ) = 1 ) then
                fin <= '0';
             end if;
          end if;
       end loop;
    end process gen_fin;

    GetCLKAPeriod : process ( CLKA_ipd, POWERDOWN_ipd, FBSEL_illegal, normalized_fb_delay, DIVN, DIVM, locked_vco0_edges, external_dly_correct )
      -- locked_vco0_edges is in the sensitivity list so that we periodically check for CLKA stopped
      variable re                 : Time :=  0.000 ns; -- Current CLKA rising edge
      variable CLKA_num_re_stable : Integer := -1;   -- Number of CLKA rising edges that PLL config stable
    begin
      if (( TO_X01( POWERDOWN_ipd ) = '1' ) and ( FBSEL_illegal = False ))  then
        if ( normalized_fb_delay'event or DIVN'event or DIVM'event or
             ( ( '1' = using_EXTFB ) and ( '1' /= external_dly_correct ) ) ) then
          internal_lock <= false;
          CLKA_num_re_stable := -1;
        end if;
        if ( CLKA_ipd'event and ( '1' = TO_X01( CLKA_ipd ) ) ) then
           if ( CLKA_period /= ( NOW - re ) ) then
              CLKA_period <= ( NOW - re );
              CLKA_num_re_stable := -1;
              internal_lock <= false;
              CLKA_period_stable <= false;
           else
              if ( f_CLKA_LOCK > CLKA_num_re_stable ) then
                 CLKA_num_re_stable := CLKA_num_re_stable + 1;
              elsif ( f_CLKA_LOCK = CLKA_num_re_stable ) then
                 internal_lock <=  true;
              end if;
              CLKA_period_stable <= true;
           end if;
           re := NOW;
        elsif ( CLKA_period < ( NOW - re ) ) then
           CLKA_num_re_stable := -1;
           internal_lock <= false;
           CLKA_period_stable <= false;
        end if;
      else
        CLKA_num_re_stable := -1;
        internal_lock <= false;
        CLKA_period_stable <= false;
      end if;
    end process GetCLKAPeriod;

    fin_period         <= CLKA_period * DIVN;

    GLA_pw             <= PLLCLK_pw * DIVU;

    extfbin_fin_drift  <= ( GLA_pw * DIVM * 2.0 ) - fin_period;

    PLLCLK_period      <= fin_period / real( fb_loop_div );

    PLLCLK_pw          <= PLLCLK_period / 2.0;

    calc_fb_loop_div : process( DIVM, DIVU, using_EXTFB )
    begin
       if ( using_EXTFB  = '1' ) then
           fb_loop_div <= DIVM * DIVU; 
       else
           fb_loop_div <= DIVM;
       end if;
    end process calc_fb_loop_div;

    sync_pll : process( fin, internal_lock, DYNSYNC )
    begin
       if ( not( internal_lock ) or ( '1' = DYNSYNC ) ) then
          locked <= '0';
       elsif ( rising_edge( fin ) ) then
          locked <= '1';
       end if;
    end process sync_pll;

    count_locked_vco0_edges: process( locked, locked_vco0_edges )
    begin
       if ( locked'event ) then
          if ( locked = '1' ) then
            locked_vco0_edges <= 0;
          else
            locked_vco0_edges <= -1;
          end if;
       elsif ( locked = '1' ) then
          if ( ( locked_vco0_edges mod( DIVU * DIVV * DIVW * DIVM * 2 ) ) = 0 ) then
             locked_vco0_edges <= 1 after PLLCLK_pw;
          else
             locked_vco0_edges <= ( locked_vco0_edges + 1 ) after PLLCLK_pw;
          end if;
       end if;
    end process count_locked_vco0_edges;

    gen_vco0_div: process( locked_vco0_edges )
    begin
       if ( locked_vco0_edges = -1 ) then
          vco0_divu <= '0';
          vco0_divv <= '0';
          vco0_divw <= '0';
       else 
         if ( ( locked_vco0_edges mod DIVU ) = 0 ) then
           vco0_divu <= not vco0_divu;
         end if;
         if ( ( locked_vco0_edges mod DIVV ) = 0 ) then
           vco0_divv <= not vco0_divv;
         end if;
         if ( ( locked_vco0_edges mod DIVW ) = 0 ) then
           vco0_divw <= not vco0_divw;
         end if;
       end if;
    end process gen_vco0_div;

    UIN <= output_mux_driver(  OAMUX_config, halveA, CLKA_ipd, CLKA2X, vco0_divu );
    VIN <= output_mux_driver(  OBMUX_config, halveB, CLKB_ipd, CLKB2X, vco0_divv );
    WIN <= output_mux_driver(  OCMUX_config, halveC, CLKC_ipd, CLKC2X, vco0_divw );

    double_CLKA: process( CLKA_ipd )
       variable re      : Time := 0 ns;
       variable prev_re : Time := 0 ns;
       variable period  : Time := 0 ns;
    begin
       if ( TO_X01( CLKA_ipd ) = '1' ) then
         prev_re := re;
         re := NOW;
         period := re - prev_re;
         if ( period > 0 ns ) then
            CLKA2X <= '1';
            CLKA2X <= transport '0' after ( period / 4.0 );
            CLKA2X <= transport '1' after ( period / 2.0 );
            CLKA2X <= transport '0' after ( period * 3.0 / 4.0 );
         end if;
       end if;
    end process double_CLKA;

    double_CLKB: process( CLKB_ipd )
       variable re      : Time := 0 ns;
       variable prev_re : Time := 0 ns;
       variable period  : Time := 0 ns;
    begin
       if ( TO_X01( CLKB_ipd ) = '1' ) then
         prev_re := re;
         re := NOW;
         period := re - prev_re;
         if ( period > 0 ns ) then
            CLKB2X <= '1';
            CLKB2X <= transport '0' after ( period / 4.0 );
            CLKB2X <= transport '1' after ( period / 2.0 );
            CLKB2X <= transport '0' after ( period * 3.0 / 4.0 );
         end if;
       end if;
    end process double_CLKB;

    double_CLKC: process( CLKC_ipd )
       variable re      : Time := 0 ns;
       variable prev_re : Time := 0 ns;
       variable period  : Time := 0 ns;
    begin
       if ( TO_X01( CLKC_ipd ) = '1' ) then
         prev_re := re;
         re := NOW;
         period := re - prev_re;
         if ( period > 0 ns ) then
            CLKC2X <= '1';
            CLKC2X <= transport '0' after ( period / 4.0 );
            CLKC2X <= transport '1' after ( period / 2.0 );
            CLKC2X <= transport '0' after ( period * 3.0 / 4.0 );
         end if;
       end if;
    end process double_CLKC;

    --
    -- AOUT Output of Divider U
    --

    DividerU : process ( UIN, CLKA_ipd, OADIVRST_ipd, OADIVHALF_ipd, 
                         POWERDOWN_ipd )

      variable force_0         : Boolean  := True;
      variable num_edges       : Integer  := -1;
      variable res_post_reset1 : Integer  :=  0;
      variable fes_post_reset1 : Integer  :=  0;
      variable res_post_reset0 : Integer  :=  0;
      variable fes_post_reset0 : Integer  :=  0;

    begin

      if ( 1 = OAMUX_config ) then -- PLL core bypassed.  OADIVRST active.

        if ( CLKA_ipd'event ) then
          if ( TO_X01( CLKA_ipd ) = '1' and TO_X01( CLKA_ipd'last_value ) = '0' ) then
             if ( 4 > res_post_reset1 ) then
                res_post_reset1 := res_post_reset1 + 1;
             end if;
             if ( 4 > res_post_reset0 ) then
               res_post_reset0 := res_post_reset0 + 1;
             end if;
             if ( res_post_reset1 = 3 ) then
                force_0 := False;
                num_edges := -1;
             end if;
          elsif ( TO_X01( CLKA_ipd ) = '0' and TO_X01( CLKA_ipd'last_value ) = '1' ) then
             if ( 4 > fes_post_reset1 ) then
               fes_post_reset1 := fes_post_reset1 + 1;
             end if;
             if ( 4 > fes_post_reset0 ) then
               fes_post_reset0 := fes_post_reset0 + 1;
             end if;
             if ( fes_post_reset1 = 1 ) then
                force_0 := True;
             end if;
          end if;
        end if;

        if ( OADIVRST_ipd'event ) then
          if ( TO_X01( OADIVRST_ipd ) = '1' ) then
            if ( ( TO_X01( OADIVRST_ipd'last_value ) = '0' ) and
                 ( ( res_post_reset0 < 1 ) or ( fes_post_reset0 < 1 ) ) ) then
              assert false
              report "OADIVRST must be held low for at least one CLKA period for the reset operation to work correctly: reset operation may not be successful, edge alignment unpredictable"
              severity warning;
            end if;
            res_post_reset1 := 0;
            fes_post_reset1 := 0;
          elsif ( TO_X01( OADIVRST_ipd ) = '0' ) then
            if ( ( TO_X01( OADIVRST_ipd'last_value ) = '1' ) and
                 ( ( res_post_reset1 < 3 ) or ( fes_post_reset1 < 3 ) ) ) then
              assert false
              report "OADIVRST must be held high for at least three CLKA periods for the reset operation to work correctly: reset operation may not be succesful, edge alignment unpredictable"
              severity warning;
            end if;
            res_post_reset0 := 0;
            fes_post_reset0 := 0;
          else
            assert false
            report "OADIVRST is unknown. Edge alignment unpredictable."
            severity warning;
          end if;
        end if;

        if ( UIN'event ) then
          num_edges := num_edges + 1;
          if ( force_0 ) then
            AOUT <= '0';
          elsif ( TO_X01( UIN ) = 'X' ) then
            AOUT <= 'X';
          elsif ( ( num_edges mod DIVU ) = 0 ) then
            num_edges := 0;
            if ( TO_X01 ( AOUT ) = 'X' ) then
              AOUT <= UIN;
            else
              AOUT <= not AOUT;
            end if;
          end if;
        end if;

      else -- PLL not bypassed
        if ( TO_X01 ( POWERDOWN_ipd ) = '0' ) then
          AOUT <= '0';
        elsif ( TO_X01 ( POWERDOWN_ipd ) = '1' ) then
          AOUT <= UIN;
        else -- POWERDOWN unknown
          AOUT <= 'X';
        end if;
      end if;

    end process DividerU;


    --
    -- BOUT Output of Divider V
    --

    DividerV : process ( VIN, CLKB_ipd, OBDIVRST_ipd, OBDIVHALF_ipd,
                         POWERDOWN_ipd )

      variable force_0         : Boolean  := True;
      variable num_edges       : Integer  := -1;
      variable res_post_reset1 : Integer  :=  0;
      variable fes_post_reset1 : Integer  :=  0;
      variable res_post_reset0 : Integer  :=  0;
      variable fes_post_reset0 : Integer  :=  0;

    begin

      if ( 0 = OBMUX_config ) then
        BOUT <= 'X';
      elsif ( 1 = OBMUX_config ) then -- PLL core bypassed.  OBDIVRST active.

        if ( CLKB_ipd'event ) then
          if ( TO_X01( CLKB_ipd ) = '1' and TO_X01( CLKB_ipd'last_value ) = '0' ) then
             if ( 4 > res_post_reset1 ) then
               res_post_reset1 := res_post_reset1 + 1;
             end if;
             if ( 4 > res_post_reset0 ) then
               res_post_reset0 := res_post_reset0 + 1;
             end if;
             if ( res_post_reset1 = 3 ) then
                force_0 := False;
                num_edges := -1;
             end if;
          elsif ( TO_X01( CLKB_ipd ) = '0' and TO_X01( CLKB_ipd'last_value ) = '1' ) then
             if ( 4 > fes_post_reset1 ) then
               fes_post_reset1 := fes_post_reset1 + 1;
             end if;
             if ( 4 > fes_post_reset0 ) then
               fes_post_reset0 := fes_post_reset0 + 1;
             end if;
             if ( fes_post_reset1 = 1 ) then
                force_0 := True;
             end if;
          end if;
        end if;

        if ( OBDIVRST_ipd'event ) then
          if ( TO_X01( OBDIVRST_ipd ) = '1' ) then
            if ( ( TO_X01( OBDIVRST_ipd'last_value ) = '0' ) and
                 ( ( res_post_reset0 < 1 ) or ( fes_post_reset0 < 1 ) ) ) then
              assert false
              report "OBDIVRST must be held low for at least one CLKB period for the reset operation to work correctly: reset operation may not be successful, edge alignment unpredictable"
              severity warning;
            end if;
            res_post_reset1 := 0;
            fes_post_reset1 := 0;
          elsif ( TO_X01( OBDIVRST_ipd ) = '0' ) then
            if ( ( TO_X01( OBDIVRST_ipd'last_value ) = '1' ) and
                 ( ( res_post_reset1 < 3 ) or ( fes_post_reset1 < 3 ) ) ) then
              assert false
              report "OBDIVRST must be held high for at least three CLKB periods for the reset operation to work correctly: reset operation may not be succesful, edge alignment unpredictable"
              severity warning;
            end if;
            res_post_reset0 := 0;
            fes_post_reset0 := 0;
          else
            assert false
            report "OBDIVRST is unknown. Edge alignment unpredictable."
            severity warning;
          end if;
        end if;

        if ( VIN'event ) then
          num_edges := num_edges + 1;
          if ( force_0 ) then
            BOUT <= '0';
          elsif ( TO_X01( VIN ) = 'X' ) then
            BOUT <= 'X';
          elsif ( ( num_edges mod DIVV ) = 0 ) then
            num_edges := 0;
            if ( TO_X01 ( BOUT ) = 'X' ) then
              BOUT <= VIN;
            else
              BOUT <= not BOUT;
            end if;
          end if;
        end if;

      else -- PLL not bypassed
        if ( TO_X01 ( POWERDOWN_ipd ) = '0' ) then
          BOUT <= '0';
        elsif ( TO_X01 ( POWERDOWN_ipd ) = '1' ) then
          BOUT <= VIN;
        else -- POWERDOWN unknown
          BOUT <= 'X';
        end if;
      end if;

    end process DividerV;

    --
    -- COUT Output of Divider W
    --

    DividerW : process ( WIN, CLKC_ipd, OCDIVRST_ipd, OCDIVHALF_ipd,
                         POWERDOWN_ipd )

      variable force_0         : Boolean  := True;
      variable num_edges       : Integer  := -1;
      variable res_post_reset1 : Integer  :=  0;
      variable fes_post_reset1 : Integer  :=  0;
      variable res_post_reset0 : Integer  :=  0;
      variable fes_post_reset0 : Integer  :=  0;

    begin

      if ( 0 = OCMUX_config ) then
        COUT <= 'X';
      elsif ( 1 = OCMUX_config ) then -- PLL core bypassed.  OCDIVRST active.

        if ( CLKC_ipd'event ) then
          if ( TO_X01( CLKC_ipd ) = '1' and TO_X01( CLKC_ipd'last_value ) = '0' ) then
             if ( 4 > res_post_reset1 ) then
               res_post_reset1 := res_post_reset1 + 1;
             end if;
             if ( 4 > res_post_reset0 ) then
               res_post_reset0 := res_post_reset0 + 1;
             end if;
             if ( res_post_reset1 = 3 ) then
                force_0 := False;
                num_edges := -1;
             end if;
          elsif ( TO_X01( CLKC_ipd ) = '0' and TO_X01( CLKC_ipd'last_value ) = '1' ) then
             if ( 4 > fes_post_reset1 ) then
               fes_post_reset1 := fes_post_reset1 + 1;
             end if;
             if ( 4 > fes_post_reset0 ) then
               fes_post_reset0 := fes_post_reset0 + 1;
             end if;
             if ( fes_post_reset1 = 1 ) then
                force_0 := True;
             end if;
          end if;
        end if;

        if ( OCDIVRST_ipd'event ) then
          if ( TO_X01( OCDIVRST_ipd ) = '1' ) then
            if ( ( TO_X01( OCDIVRST_ipd'last_value ) = '0' ) and
                 ( ( res_post_reset0 < 1 ) or ( fes_post_reset0 < 1 ) ) ) then
              assert false
              report "OCDIVRST must be held low for at least one CLKC period for the reset operation to work correctly: reset operation may not be successful, edge alignment unpredictable"
              severity warning;
            end if;
            res_post_reset1 := 0;
            fes_post_reset1 := 0;
          elsif ( TO_X01( OCDIVRST_ipd ) = '0' ) then
            if ( ( TO_X01( OCDIVRST_ipd'last_value ) = '1' ) and
                 ( ( res_post_reset1 < 3 ) or ( fes_post_reset1 < 3 ) ) ) then
              assert false
              report "OCDIVRST must be held high for at least three CLKC periods for the reset operation to work correctly: reset operation may not be succesful, edge alignment unpredictable"
              severity warning;
            end if;
            res_post_reset0 := 0;
            fes_post_reset0 := 0;
          else
            assert false
            report "OCDIVRST is unknown. Edge alignment unpredictable."
            severity warning;
          end if;
        end if;

        if ( WIN'event ) then
          num_edges := num_edges + 1;
          if ( force_0 ) then
            COUT <= '0';
          elsif ( TO_X01( WIN ) = 'X' ) then
            COUT <= 'X';
          elsif ( ( num_edges mod DIVW ) = 0 ) then
            num_edges := 0;
            if ( TO_X01 ( COUT ) = 'X' ) then
              COUT <= WIN;
            else
              COUT <= not COUT;
            end if;
          end if;
        end if;

      else -- PLL not bypassed
        if ( TO_X01 ( POWERDOWN_ipd ) = '0' ) then
          COUT <= '0';
        elsif ( TO_X01 ( POWERDOWN_ipd ) = '1' ) then
          COUT <= WIN;
        else -- POWERDOWN unknown
          COUT <= 'X';
        end if;
      end if;

    end process DividerW;

    using_EXTFB <= TO_X01( FBSEL1_ipd and FBSEL0_ipd );

    external_dly_correct <= expected_EXTFB xnor EXTFB_ipd after 1 ps;

    get_EXTFB_period : process
      variable previous_re : time :=  0.000 ns; -- Previous EXTFB rising edge
    begin
      wait until rising_edge( EXTFB );
      EXTFB_period <= NOW - previous_re;
      previous_re := NOW;
    end process get_EXTFB_period;

    calculate_extfb_delay : process
      variable CLKA_edge : time := 0 ns;
    begin
       EXTFB_delay_dtrmd <= false;
       if ( ( '1' /= using_EXTFB ) or ( not CLKA_period_stable ) ) then
          wait until ( ( '1' = using_EXTFB ) and CLKA_period_stable );
       end if;
       wait for GLA_EXTFB_rise_dly;
       GLA_EXTFB_fall_dly <= 0 ps;
       GLA_EXTFB_rise_dly <= 0 ps;
       wait for ( CLKA_2_GLA_dly * 2);
       calibrate_EXTFB_delay <= '1';
       if ( '1' /= EXTFB_ipd ) then
          wait until ( EXTFB_ipd = '1' );
       end if;
       wait until falling_edge( CLKA_ipd );
       CLKA_edge := NOW;
       calibrate_EXTFB_delay <= '0';
       wait until falling_edge( EXTFB_ipd );
       GLA_EXTFB_fall_dly <= NOW - CLKA_edge - CLKA_2_GLA_dly;
       wait until rising_edge( CLKA_ipd );
       CLKA_edge := NOW;
       calibrate_EXTFB_delay <= '1';
       wait until rising_edge( EXTFB_ipd );
       GLA_EXTFB_rise_dly <= NOW - CLKA_edge - CLKA_2_GLA_dly;
       wait until falling_edge( CLKA_ipd );
       wait until ( CLKA_period_stable and rising_edge( fin ) );
       EXTFB_delay_dtrmd <= true;
       wait until falling_edge( expected_EXTFB );
       if ( '1' /= external_dly_correct ) then
         assert false
         report "ERROR: EXTFB must be a simple, time-delayed derivative of GLA. Simulation cannot continue until user-logic is corrected"
         severity failure;
         wait;
       end if;
       wait until ( '1' /= external_dly_correct );
    end process calculate_extfb_delay;

    external_feedback : process
       variable edges : integer := 1;
    begin
       wait on GLA_free_running, EXTFB_delay_dtrmd;
       if ( EXTFB_delay_dtrmd ) then
         if ( ( edges mod ( DIVM * 2 ) ) = 0 ) then
            GLA_free_running <= not GLA_free_running after ( GLA_pw - extfbin_fin_drift );
            edges := 0;
         else
            GLA_free_running <= not GLA_free_running after GLA_pw;
         end if;
         edges := edges + 1;
       else
         edges := 1;
         GLA_free_running <= '1' after GLA_pw;
       end if;
    end process external_feedback;

    gen_AOUT_using_EXTFB : process( AOUT, GLA_free_running, calibrate_EXTFB_delay, locked_vco0_edges, EXTFB_delay_dtrmd )
    begin
       if ( 0 <= locked_vco0_edges ) then
          AOUT_using_EXTFB <= AOUT;
       elsif ( EXTFB_delay_dtrmd ) then
          AOUT_using_EXTFB <= GLA_free_running;
       else
          AOUT_using_EXTFB <= calibrate_EXTFB_delay;
       end if;
    end process gen_AOUT_using_EXTFB;

    gen_expected_EXTFB: process( AOUT_using_EXTFB, EXTFB_delay_dtrmd )
    begin
       if ( not EXTFB_delay_dtrmd ) then
          expected_EXTFB <= 'X';
       elsif ( '1' = AOUT_using_EXTFB ) then
          expected_EXTFB <= transport AOUT_using_EXTFB after ( CLKA_2_GLA_dly + GLA_EXTFB_rise_dly );
       else
          expected_EXTFB <= transport AOUT_using_EXTFB after ( CLKA_2_GLA_dly + GLA_EXTFB_fall_dly );
       end if;
    end process gen_expected_EXTFB;

    Aoutputs: process( AOUT, CLKA_ipd, AOUT_using_EXTFB, OAMUX_config  )
    begin
        if ( 0 = OAMUX_config ) then
          GLA <= transport CLKA_ipd after CLKA_2_GLA_bypass0_dly;
        elsif ( ( 1 = OAMUX_config ) or ( 3 = OAMUX_config ) ) then
          GLA <= transport 'X' after CLKA_2_GLA_dly;
          assert ( not OAMUX_config'event )
            report "WARNING: Illegal OAMUX configuration."
            severity warning;
        elsif ( '1' = using_EXTFB ) then
          GLA <= transport AOUT_using_EXTFB after CLKA_2_GLA_dly;
        else
          GLA <= transport AOUT after CLKA_2_GLA_dly;
        end if;
    end process Aoutputs;
    
    Boutputs: process ( BOUT, CLKB_ipd, OBMUX_config )
    begin
        if ( 0 = OBMUX_config ) then
          GLB <= transport CLKB_ipd after CLKB_2_GLB_bypass0_dly;
          YB  <= 'X';
        elsif ( ( 1 = OBMUX_config ) or ( 3 = OBMUX_config ) ) then
          GLB <= transport 'X' after CLKA_2_GLB_dly;
          YB  <= transport 'X' after CLKA_2_YB_dly;
          assert ( not OBMUX_config'event )
            report "WARNING: Illegal OBMUX configuration."
            severity warning;
        else
          GLB <= transport BOUT after CLKA_2_GLB_dly;
          YB  <= transport BOUT after CLKA_2_YB_dly;
        end if;
    end process Boutputs;

    Coutputs: process ( COUT, CLKC_ipd, OCMUX_config )
    begin
        if ( 0 = OCMUX_config ) then
          GLC <= transport CLKC_ipd after CLKC_2_GLC_bypass0_dly;
          YC  <= 'X';
        elsif ( ( 1 = OCMUX_config ) or ( 3 = OCMUX_config ) ) then
          GLC <= transport 'X' after CLKA_2_GLC_dly;
          YC  <= transport 'X' after CLKA_2_YC_dly;
          assert ( not OCMUX_config'event )
            report "WARNING: Illegal OCMUX configuration."
            severity warning;
        else
          GLC <= transport COUT after CLKA_2_GLC_dly;
          YC  <= transport COUT after CLKA_2_YC_dly;
        end if;
    end process Coutputs;
    
  end VITAL_ACT;

configuration CFG_PLLPRIM_VITAL of PLLPRIM is
  for VITAL_ACT
  end for;
end CFG_PLLPRIM_VITAL;

----- CELL PLL -----

library IEEE;
use IEEE.std_logic_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
 entity PLL is
  generic(
    VCOFREQUENCY      :  Real    := 0.0;
    f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

    TimingChecksOn    :  Boolean          := True;
    InstancePath      :  String           := "*";
    Xon               :  Boolean          := False;
    MsgOn             :  Boolean          := True;
    
    tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV5      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV6      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV5       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV6       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBSEL0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBSEL1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_XDLYSEL      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

    tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns )
   );

  port (
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    POWERDOWN    : in    std_ulogic;
    OADIV0       : in    std_ulogic;
    OADIV1       : in    std_ulogic;
    OADIV2       : in    std_ulogic;
    OADIV3       : in    std_ulogic;
    OADIV4       : in    std_ulogic;
    OAMUX0       : in    std_ulogic;
    OAMUX1       : in    std_ulogic;
    OAMUX2       : in    std_ulogic;
    DLYGLA0      : in    std_ulogic;
    DLYGLA1      : in    std_ulogic;
    DLYGLA2      : in    std_ulogic;
    DLYGLA3      : in    std_ulogic;
    DLYGLA4      : in    std_ulogic;
    OBDIV0       : in    std_ulogic;
    OBDIV1       : in    std_ulogic;
    OBDIV2       : in    std_ulogic;
    OBDIV3       : in    std_ulogic;
    OBDIV4       : in    std_ulogic;
    OBMUX0       : in    std_ulogic;
    OBMUX1       : in    std_ulogic;
    OBMUX2       : in    std_ulogic;
    DLYYB0       : in    std_ulogic;
    DLYYB1       : in    std_ulogic;
    DLYYB2       : in    std_ulogic;
    DLYYB3       : in    std_ulogic;
    DLYYB4       : in    std_ulogic;
    DLYGLB0      : in    std_ulogic;
    DLYGLB1      : in    std_ulogic;
    DLYGLB2      : in    std_ulogic;
    DLYGLB3      : in    std_ulogic;
    DLYGLB4      : in    std_ulogic;
    OCDIV0       : in    std_ulogic;
    OCDIV1       : in    std_ulogic;
    OCDIV2       : in    std_ulogic;
    OCDIV3       : in    std_ulogic;
    OCDIV4       : in    std_ulogic;
    OCMUX0       : in    std_ulogic;
    OCMUX1       : in    std_ulogic;
    OCMUX2       : in    std_ulogic;
    DLYYC0       : in    std_ulogic;
    DLYYC1       : in    std_ulogic;
    DLYYC2       : in    std_ulogic;
    DLYYC3       : in    std_ulogic;
    DLYYC4       : in    std_ulogic;
    DLYGLC0      : in    std_ulogic;
    DLYGLC1      : in    std_ulogic;
    DLYGLC2      : in    std_ulogic;
    DLYGLC3      : in    std_ulogic;
    DLYGLC4      : in    std_ulogic;
    FINDIV0      : in    std_ulogic;
    FINDIV1      : in    std_ulogic;
    FINDIV2      : in    std_ulogic;
    FINDIV3      : in    std_ulogic;
    FINDIV4      : in    std_ulogic;
    FINDIV5      : in    std_ulogic;
    FINDIV6      : in    std_ulogic;
    FBDIV0       : in    std_ulogic;
    FBDIV1       : in    std_ulogic;
    FBDIV2       : in    std_ulogic;
    FBDIV3       : in    std_ulogic;
    FBDIV4       : in    std_ulogic;
    FBDIV5       : in    std_ulogic;
    FBDIV6       : in    std_ulogic;
    FBDLY0       : in    std_ulogic;
    FBDlY1       : in    std_ulogic;
    FBDLY2       : in    std_ulogic;
    FBDLY3       : in    std_ulogic;
    FBDlY4       : in    std_ulogic;
    FBSEL0       : in    std_ulogic;
    FBSEL1       : in    std_ulogic;
    XDLYSEL      : in    std_ulogic;
    VCOSEL0      : in    std_ulogic;
    VCOSEL1      : in    std_ulogic;
    VCOSEL2      : in    std_ulogic;
    GLA          : out   std_ulogic;
    LOCK         : out   std_ulogic;
    GLB          : out   std_ulogic;
    YB           : out   std_ulogic;
    GLC          : out   std_ulogic;
    YC           : out   std_ulogic
   );

  attribute VITAL_LEVEL0 of PLL : entity is TRUE;
end PLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.components.all;

architecture VITAL_ACT of PLL is
attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal CLKA_ipd               : std_ulogic;
  signal EXTFB_ipd              : std_ulogic;
  signal POWERDOWN_ipd          : std_ulogic;
  signal OADIV0_ipd             : std_ulogic;
  signal OADIV1_ipd             : std_ulogic;
  signal OADIV2_ipd             : std_ulogic;
  signal OADIV3_ipd             : std_ulogic;
  signal OADIV4_ipd             : std_ulogic;
  signal OAMUX0_ipd             : std_ulogic;
  signal OAMUX1_ipd             : std_ulogic;
  signal OAMUX2_ipd             : std_ulogic;
  signal DLYGLA0_ipd            : std_ulogic;
  signal DLYGLA1_ipd            : std_ulogic;
  signal DLYGLA2_ipd            : std_ulogic;
  signal DLYGLA3_ipd            : std_ulogic;
  signal DLYGLA4_ipd            : std_ulogic;
  signal OBDIV0_ipd             : std_ulogic;
  signal OBDIV1_ipd             : std_ulogic;
  signal OBDIV2_ipd             : std_ulogic;
  signal OBDIV3_ipd             : std_ulogic;
  signal OBDIV4_ipd             : std_ulogic;
  signal OBMUX0_ipd             : std_ulogic;
  signal OBMUX1_ipd             : std_ulogic;
  signal OBMUX2_ipd             : std_ulogic;
  signal DLYYB0_ipd             : std_ulogic;
  signal DLYYB1_ipd             : std_ulogic;
  signal DLYYB2_ipd             : std_ulogic;
  signal DLYYB3_ipd             : std_ulogic;
  signal DLYYB4_ipd             : std_ulogic;
  signal DLYGLB0_ipd            : std_ulogic;
  signal DLYGLB1_ipd            : std_ulogic;
  signal DLYGLB2_ipd            : std_ulogic;
  signal DLYGLB3_ipd            : std_ulogic;
  signal DLYGLB4_ipd            : std_ulogic;
  signal OCDIV0_ipd             : std_ulogic;
  signal OCDIV1_ipd             : std_ulogic;
  signal OCDIV2_ipd             : std_ulogic;
  signal OCDIV3_ipd             : std_ulogic;
  signal OCDIV4_ipd             : std_ulogic;
  signal OCMUX0_ipd             : std_ulogic;
  signal OCMUX1_ipd             : std_ulogic;
  signal OCMUX2_ipd             : std_ulogic;
  signal DLYYC0_ipd             : std_ulogic;
  signal DLYYC1_ipd             : std_ulogic;
  signal DLYYC2_ipd             : std_ulogic;
  signal DLYYC3_ipd             : std_ulogic;
  signal DLYYC4_ipd             : std_ulogic;
  signal DLYGLC0_ipd            : std_ulogic;
  signal DLYGLC1_ipd            : std_ulogic;
  signal DLYGLC2_ipd            : std_ulogic;
  signal DLYGLC3_ipd            : std_ulogic;
  signal DLYGLC4_ipd            : std_ulogic;
  signal FINDIV0_ipd            : std_ulogic;
  signal FINDIV1_ipd            : std_ulogic;
  signal FINDIV2_ipd            : std_ulogic;
  signal FINDIV3_ipd            : std_ulogic;
  signal FINDIV4_ipd            : std_ulogic;
  signal FINDIV5_ipd            : std_ulogic;
  signal FINDIV6_ipd            : std_ulogic;
  signal FBDIV0_ipd             : std_ulogic;
  signal FBDIV1_ipd             : std_ulogic;
  signal FBDIV2_ipd             : std_ulogic;
  signal FBDIV3_ipd             : std_ulogic;
  signal FBDIV4_ipd             : std_ulogic;
  signal FBDIV5_ipd             : std_ulogic;
  signal FBDIV6_ipd             : std_ulogic;
  signal FBDLY0_ipd             : std_ulogic;
  signal FBDlY1_ipd             : std_ulogic;
  signal FBDLY2_ipd             : std_ulogic;
  signal FBDLY3_ipd             : std_ulogic;
  signal FBDlY4_ipd             : std_ulogic;
  signal FBSEL0_ipd             : std_ulogic;
  signal FBSEL1_ipd             : std_ulogic;
  signal XDLYSEL_ipd            : std_ulogic;
  signal VCOSEL0_ipd            : std_ulogic;
  signal VCOSEL1_ipd            : std_ulogic;
  signal VCOSEL2_ipd            : std_ulogic;

  signal GND                    : std_logic := '0';
  signal UNUSED                 : std_logic := 'X';

  component PLLPRIM
    generic (
              VCOFREQUENCY :  Real;
              f_CLKA_LOCK  :  Integer
            );
    port (
           DYNSYNC      : in    std_ulogic;
           CLKA         : in    std_ulogic;
           EXTFB        : in    std_ulogic;
           POWERDOWN    : in    std_ulogic;
           CLKB         : in    std_ulogic;
           CLKC         : in    std_ulogic;
           OADIVRST     : in    std_ulogic;
           OADIVHALF    : in    std_ulogic;
           OADIV0       : in    std_ulogic;
           OADIV1       : in    std_ulogic;
           OADIV2       : in    std_ulogic;
           OADIV3       : in    std_ulogic;
           OADIV4       : in    std_ulogic;
           OAMUX0       : in    std_ulogic;
           OAMUX1       : in    std_ulogic;
           OAMUX2       : in    std_ulogic;
           DLYGLA0      : in    std_ulogic;
           DLYGLA1      : in    std_ulogic;
           DLYGLA2      : in    std_ulogic;
           DLYGLA3      : in    std_ulogic;
           DLYGLA4      : in    std_ulogic;
           OBDIVRST     : in    std_ulogic;
           OBDIVHALF    : in    std_ulogic;
           OBDIV0       : in    std_ulogic;
           OBDIV1       : in    std_ulogic;
           OBDIV2       : in    std_ulogic;
           OBDIV3       : in    std_ulogic;
           OBDIV4       : in    std_ulogic;
           OBMUX0       : in    std_ulogic;
           OBMUX1       : in    std_ulogic;
           OBMUX2       : in    std_ulogic;
           DLYYB0       : in    std_ulogic;
           DLYYB1       : in    std_ulogic;
           DLYYB2       : in    std_ulogic;
           DLYYB3       : in    std_ulogic;
           DLYYB4       : in    std_ulogic;
           DLYGLB0      : in    std_ulogic;
           DLYGLB1      : in    std_ulogic;
           DLYGLB2      : in    std_ulogic;
           DLYGLB3      : in    std_ulogic;
           DLYGLB4      : in    std_ulogic;
           OCDIVRST     : in    std_ulogic;
           OCDIVHALF    : in    std_ulogic;
           OCDIV0       : in    std_ulogic;
           OCDIV1       : in    std_ulogic;
           OCDIV2       : in    std_ulogic;
           OCDIV3       : in    std_ulogic;
           OCDIV4       : in    std_ulogic;
           OCMUX0       : in    std_ulogic;
           OCMUX1       : in    std_ulogic;
           OCMUX2       : in    std_ulogic;
           DLYYC0       : in    std_ulogic;
           DLYYC1       : in    std_ulogic;
           DLYYC2       : in    std_ulogic;
           DLYYC3       : in    std_ulogic;
           DLYYC4       : in    std_ulogic;
           DLYGLC0      : in    std_ulogic;
           DLYGLC1      : in    std_ulogic;
           DLYGLC2      : in    std_ulogic;
           DLYGLC3      : in    std_ulogic;
           DLYGLC4      : in    std_ulogic;
           FINDIV0      : in    std_ulogic;
           FINDIV1      : in    std_ulogic;
           FINDIV2      : in    std_ulogic;
           FINDIV3      : in    std_ulogic;
           FINDIV4      : in    std_ulogic;
           FINDIV5      : in    std_ulogic;
           FINDIV6      : in    std_ulogic;
           FBDIV0       : in    std_ulogic;
           FBDIV1       : in    std_ulogic;
           FBDIV2       : in    std_ulogic;
           FBDIV3       : in    std_ulogic;
           FBDIV4       : in    std_ulogic;
           FBDIV5       : in    std_ulogic;
           FBDIV6       : in    std_ulogic;
           FBDLY0       : in    std_ulogic;
           FBDlY1       : in    std_ulogic;
           FBDLY2       : in    std_ulogic;
           FBDLY3       : in    std_ulogic;
           FBDlY4       : in    std_ulogic;
           FBSEL0       : in    std_ulogic;
           FBSEL1       : in    std_ulogic;
           XDLYSEL      : in    std_ulogic;
           VCOSEL0      : in    std_ulogic;
           VCOSEL1      : in    std_ulogic;
           VCOSEL2      : in    std_ulogic;
           GLA          : out   std_ulogic;
           LOCK         : out   std_ulogic;
           GLB          : out   std_ulogic;
           YB           : out   std_ulogic;
           GLC          : out   std_ulogic;
           YC           : out   std_ulogic
         );
  end component;

  begin

    ---------------------
    --  INPUT PATH DELAYs
    ---------------------
    WireDelay : block

    begin

      VitalWireDelay ( CLKA_ipd,      CLKA,      tipd_CLKA );
      VitalWireDelay ( EXTFB_ipd,     EXTFB,     tipd_EXTFB );
      VitalWireDelay ( POWERDOWN_ipd, POWERDOWN, tipd_POWERDOWN );
      VitalWireDelay ( OADIV0_ipd,    OADIV0,    tipd_OADIV0 );
      VitalWireDelay ( OADIV1_ipd,    OADIV1,    tipd_OADIV1 );
      VitalWireDelay ( OADIV2_ipd,    OADIV2,    tipd_OADIV2 );
      VitalWireDelay ( OADIV3_ipd,    OADIV3,    tipd_OADIV3 );
      VitalWireDelay ( OADIV4_ipd,    OADIV4,    tipd_OADIV4 );
      VitalWireDelay ( OAMUX0_ipd,    OAMUX0,    tipd_OAMUX0 );
      VitalWireDelay ( OAMUX1_ipd,    OAMUX1,    tipd_OAMUX1 );
      VitalWireDelay ( OAMUX2_ipd,    OAMUX2,    tipd_OAMUX2 );
      VitalWireDelay ( DLYGLA0_ipd,   DLYGLA0,   tipd_DLYGLA0 );
      VitalWireDelay ( DLYGLA1_ipd,   DLYGLA1,   tipd_DLYGLA1 );
      VitalWireDelay ( DLYGLA2_ipd,   DLYGLA2,   tipd_DLYGLA2 );
      VitalWireDelay ( DLYGLA3_ipd,   DLYGLA3,   tipd_DLYGLA3 );
      VitalWireDelay ( DLYGLA4_ipd,   DLYGLA4,   tipd_DLYGLA4 );
      VitalWireDelay ( OBDIV0_ipd,    OBDIV0,    tipd_OBDIV0 );
      VitalWireDelay ( OBDIV1_ipd,    OBDIV1,    tipd_OBDIV1 );
      VitalWireDelay ( OBDIV2_ipd,    OBDIV2,    tipd_OBDIV2 );
      VitalWireDelay ( OBDIV3_ipd,    OBDIV3,    tipd_OBDIV3 );
      VitalWireDelay ( OBDIV4_ipd,    OBDIV4,    tipd_OBDIV4 );
      VitalWireDelay ( OBMUX0_ipd,    OBMUX0,    tipd_OBMUX0 );
      VitalWireDelay ( OBMUX1_ipd,    OBMUX1,    tipd_OBMUX1 );
      VitalWireDelay ( OBMUX2_ipd,    OBMUX2,    tipd_OBMUX2 );
      VitalWireDelay ( DLYYB0_ipd,    DLYYB0,    tipd_DLYYB0 );
      VitalWireDelay ( DLYYB1_ipd,    DLYYB1,    tipd_DLYYB1 );
      VitalWireDelay ( DLYYB2_ipd,    DLYYB2,    tipd_DLYYB2 );
      VitalWireDelay ( DLYYB3_ipd,    DLYYB3,    tipd_DLYYB3 );
      VitalWireDelay ( DLYYB4_ipd,    DLYYB4,    tipd_DLYYB4 );
      VitalWireDelay ( DLYGLB0_ipd,   DLYGLB0,   tipd_DLYGLB0 );
      VitalWireDelay ( DLYGLB1_ipd,   DLYGLB1,   tipd_DLYGLB1 );
      VitalWireDelay ( DLYGLB2_ipd,   DLYGLB2,   tipd_DLYGLB2 );
      VitalWireDelay ( DLYGLB3_ipd,   DLYGLB3,   tipd_DLYGLB3 );
      VitalWireDelay ( DLYGLB4_ipd,   DLYGLB4,   tipd_DLYGLB4 );
      VitalWireDelay ( OCDIV0_ipd,    OCDIV0,    tipd_OCDIV0 );
      VitalWireDelay ( OCDIV1_ipd,    OCDIV1,    tipd_OCDIV1 );
      VitalWireDelay ( OCDIV2_ipd,    OCDIV2,    tipd_OCDIV2 );
      VitalWireDelay ( OCDIV3_ipd,    OCDIV3,    tipd_OCDIV3 );
      VitalWireDelay ( OCDIV4_ipd,    OCDIV4,    tipd_OCDIV4 );
      VitalWireDelay ( OCMUX0_ipd,    OCMUX0,    tipd_OCMUX0 );
      VitalWireDelay ( OCMUX1_ipd,    OCMUX1,    tipd_OCMUX1 );
      VitalWireDelay ( OCMUX2_ipd,    OCMUX2,    tipd_OCMUX2 );
      VitalWireDelay ( DLYYC0_ipd,    DLYYC0,    tipd_DLYYC0 );
      VitalWireDelay ( DLYYC1_ipd,    DLYYC1,    tipd_DLYYC1 );
      VitalWireDelay ( DLYYC2_ipd,    DLYYC2,    tipd_DLYYC2 );
      VitalWireDelay ( DLYYC3_ipd,    DLYYC3,    tipd_DLYYC3 );
      VitalWireDelay ( DLYYC4_ipd,    DLYYC4,    tipd_DLYYC4 );
      VitalWireDelay ( DLYGLC0_ipd,   DLYGLC0,   tipd_DLYGLC0 );
      VitalWireDelay ( DLYGLC1_ipd,   DLYGLC1,   tipd_DLYGLC1 );
      VitalWireDelay ( DLYGLC2_ipd,   DLYGLC2,   tipd_DLYGLC2 );
      VitalWireDelay ( DLYGLC3_ipd,   DLYGLC3,   tipd_DLYGLC3 );
      VitalWireDelay ( DLYGLC4_ipd,   DLYGLC4,   tipd_DLYGLC4 );
      VitalWireDelay ( FINDIV0_ipd,   FINDIV0,   tipd_FINDIV0 );
      VitalWireDelay ( FINDIV1_ipd,   FINDIV1,   tipd_FINDIV1 );
      VitalWireDelay ( FINDIV2_ipd,   FINDIV2,   tipd_FINDIV2 );
      VitalWireDelay ( FINDIV3_ipd,   FINDIV3,   tipd_FINDIV3 );
      VitalWireDelay ( FINDIV4_ipd,   FINDIV4,   tipd_FINDIV4 );
      VitalWireDelay ( FINDIV5_ipd,   FINDIV5,   tipd_FINDIV5 );
      VitalWireDelay ( FINDIV6_ipd,   FINDIV6,   tipd_FINDIV6 );
      VitalWireDelay ( FBDIV0_ipd,    FBDIV0,    tipd_FBDIV0 );
      VitalWireDelay ( FBDIV1_ipd,    FBDIV1,    tipd_FBDIV1 );
      VitalWireDelay ( FBDIV2_ipd,    FBDIV2,    tipd_FBDIV2 );
      VitalWireDelay ( FBDIV3_ipd,    FBDIV3,    tipd_FBDIV3 );
      VitalWireDelay ( FBDIV4_ipd,    FBDIV4,    tipd_FBDIV4 );
      VitalWireDelay ( FBDIV5_ipd,    FBDIV5,    tipd_FBDIV5 );
      VitalWireDelay ( FBDIV6_ipd,    FBDIV6,    tipd_FBDIV6 );
      VitalWireDelay ( FBDLY0_ipd,    FBDLY0,    tipd_FBDLY0 );
      VitalWireDelay ( FBDLY1_ipd,    FBDLY1,    tipd_FBDLY1 );
      VitalWireDelay ( FBDLY2_ipd,    FBDLY2,    tipd_FBDLY2 );
      VitalWireDelay ( FBDLY3_ipd,    FBDLY3,    tipd_FBDLY3 );
      VitalWireDelay ( FBDLY4_ipd,    FBDLY4,    tipd_FBDLY4 );
      VitalWireDelay ( FBSEL0_ipd,    FBSEL0,    tipd_FBSEL0 );
      VitalWireDelay ( FBSEL1_ipd,    FBSEL1,    tipd_FBSEL1 );
      VitalWireDelay ( XDLYSEL_ipd,   XDLYSEL,   tipd_XDLYSEL );
      VitalWireDelay ( VCOSEL0_ipd,   VCOSEL0,   tipd_VCOSEL0 );
      VitalWireDelay ( VCOSEL1_ipd,   VCOSEL1,   tipd_VCOSEL1 );
      VitalWireDelay ( VCOSEL2_ipd,   VCOSEL2,   tipd_VCOSEL2 );
 
    end block WireDelay;
    
    P1: PLLPRIM
          generic map (
                        VCOFREQUENCY => VCOFREQUENCY,
                        f_CLKA_LOCK  => f_CLKA_LOCK
                      )
          port map    (
                        DYNSYNC      => GND,
                        CLKA         => CLKA_ipd,
                        EXTFB        => EXTFB_ipd,
                        POWERDOWN    => POWERDOWN_ipd,
                        CLKB         => UNUSED,
                        CLKC         => UNUSED,
                        OADIVRST     => GND,
                        OADIVHALF    => GND,
                        OADIV0       => OADIV0_ipd,
                        OADIV1       => OADIV1_ipd,
                        OADIV2       => OADIV2_ipd,
                        OADIV3       => OADIV3_ipd,
                        OADIV4       => OADIV4_ipd,
                        OAMUX0       => OAMUX0_ipd,
                        OAMUX1       => OAMUX1_ipd,
                        OAMUX2       => OAMUX2_ipd,
                        DLYGLA0      => DLYGLA0_ipd,
                        DLYGLA1      => DLYGLA1_ipd,
                        DLYGLA2      => DLYGLA2_ipd,
                        DLYGLA3      => DLYGLA3_ipd,
                        DLYGLA4      => DLYGLA4_ipd,
                        OBDIVRST     => GND,
                        OBDIVHALF    => GND,
                        OBDIV0       => OBDIV0_ipd,
                        OBDIV1       => OBDIV1_ipd,
                        OBDIV2       => OBDIV2_ipd,
                        OBDIV3       => OBDIV3_ipd,
                        OBDIV4       => OBDIV4_ipd,
                        OBMUX0       => OBMUX0_ipd,
                        OBMUX1       => OBMUX1_ipd,
                        OBMUX2       => OBMUX2_ipd,
                        DLYYB0       => DLYYB0_ipd,
                        DLYYB1       => DLYYB1_ipd,
                        DLYYB2       => DLYYB2_ipd,
                        DLYYB3       => DLYYB3_ipd,
                        DLYYB4       => DLYYB4_ipd,
                        DLYGLB0      => DLYGLB0_ipd,
                        DLYGLB1      => DLYGLB1_ipd,
                        DLYGLB2      => DLYGLB2_ipd,
                        DLYGLB3      => DLYGLB3_ipd,
                        DLYGLB4      => DLYGLB4_ipd,
                        OCDIVRST     => GND,
                        OCDIVHALF    => GND,
                        OCDIV0       => OCDIV0_ipd,
                        OCDIV1       => OCDIV1_ipd,
                        OCDIV2       => OCDIV2_ipd,
                        OCDIV3       => OCDIV3_ipd,
                        OCDIV4       => OCDIV4_ipd,
                        OCMUX0       => OCMUX0_ipd,
                        OCMUX1       => OCMUX1_ipd,
                        OCMUX2       => OCMUX2_ipd,
                        DLYYC0       => DLYYC0_ipd,
                        DLYYC1       => DLYYC1_ipd,
                        DLYYC2       => DLYYC2_ipd,
                        DLYYC3       => DLYYC3_ipd,
                        DLYYC4       => DLYYC4_ipd,
                        DLYGLC0      => DLYGLC0_ipd,
                        DLYGLC1      => DLYGLC1_ipd,
                        DLYGLC2      => DLYGLC2_ipd,
                        DLYGLC3      => DLYGLC3_ipd,
                        DLYGLC4      => DLYGLC4_ipd,
                        FINDIV0      => FINDIV0_ipd,
                        FINDIV1      => FINDIV1_ipd,
                        FINDIV2      => FINDIV2_ipd,
                        FINDIV3      => FINDIV3_ipd,
                        FINDIV4      => FINDIV4_ipd,
                        FINDIV5      => FINDIV5_ipd,
                        FINDIV6      => FINDIV6_ipd,
                        FBDIV0       => FBDIV0_ipd,
                        FBDIV1       => FBDIV1_ipd,
                        FBDIV2       => FBDIV2_ipd,
                        FBDIV3       => FBDIV3_ipd,
                        FBDIV4       => FBDIV4_ipd,
                        FBDIV5       => FBDIV5_ipd,
                        FBDIV6       => FBDIV6_ipd,
                        FBDLY0       => FBDLY0_ipd,
                        FBDlY1       => FBDlY1_ipd,
                        FBDLY2       => FBDLY2_ipd,
                        FBDLY3       => FBDLY3_ipd,
                        FBDlY4       => FBDlY4_ipd,
                        FBSEL0       => FBSEL0_ipd,
                        FBSEL1       => FBSEL1_ipd,
                        XDLYSEL      => XDLYSEL_ipd,
                        VCOSEL0      => VCOSEL0_ipd,
                        VCOSEL1      => VCOSEL1_ipd,
                        VCOSEL2      => VCOSEL2_ipd,
                        GLA          => GLA,
                        LOCK         => LOCK,
                        GLB          => GLB,
                        YB           => YB,
                        GLC          => GLC,
                        YC           => YC
                      );
  end VITAL_ACT;

configuration CFG_PLL_VITAL of PLL is
  for VITAL_ACT
  end for;
end CFG_PLL_VITAL;

----- CELL PLL_V2 -----

library IEEE;
use IEEE.std_logic_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
 entity PLL_V2 is
  generic(
    VCOFREQUENCY      :  Real    := 0.0;
    f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

    TimingChecksOn    :  Boolean          := True;
    InstancePath      :  String           := "*";
    Xon               :  Boolean          := False;
    MsgOn             :  Boolean          := True;
    
    tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OADIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OAMUX2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLA4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OBMUX2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYB4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLB4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_OCMUX2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYYC4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_DLYGLC4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV3      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV4      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV5      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FINDIV6      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV5       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDIV6       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY2       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY3       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBDLY4       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBSEL0       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_FBSEL1       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_XDLYSEL      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL0      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL1      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_VCOSEL2      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

    tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
    tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns )
   );

  port (
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    POWERDOWN    : in    std_ulogic;
    OADIV0       : in    std_ulogic;
    OADIV1       : in    std_ulogic;
    OADIV2       : in    std_ulogic;
    OADIV3       : in    std_ulogic;
    OADIV4       : in    std_ulogic;
    OAMUX0       : in    std_ulogic;
    OAMUX1       : in    std_ulogic;
    OAMUX2       : in    std_ulogic;
    DLYGLA0      : in    std_ulogic;
    DLYGLA1      : in    std_ulogic;
    DLYGLA2      : in    std_ulogic;
    DLYGLA3      : in    std_ulogic;
    DLYGLA4      : in    std_ulogic;
    OBDIV0       : in    std_ulogic;
    OBDIV1       : in    std_ulogic;
    OBDIV2       : in    std_ulogic;
    OBDIV3       : in    std_ulogic;
    OBDIV4       : in    std_ulogic;
    OBMUX0       : in    std_ulogic;
    OBMUX1       : in    std_ulogic;
    OBMUX2       : in    std_ulogic;
    DLYYB0       : in    std_ulogic;
    DLYYB1       : in    std_ulogic;
    DLYYB2       : in    std_ulogic;
    DLYYB3       : in    std_ulogic;
    DLYYB4       : in    std_ulogic;
    DLYGLB0      : in    std_ulogic;
    DLYGLB1      : in    std_ulogic;
    DLYGLB2      : in    std_ulogic;
    DLYGLB3      : in    std_ulogic;
    DLYGLB4      : in    std_ulogic;
    OCDIV0       : in    std_ulogic;
    OCDIV1       : in    std_ulogic;
    OCDIV2       : in    std_ulogic;
    OCDIV3       : in    std_ulogic;
    OCDIV4       : in    std_ulogic;
    OCMUX0       : in    std_ulogic;
    OCMUX1       : in    std_ulogic;
    OCMUX2       : in    std_ulogic;
    DLYYC0       : in    std_ulogic;
    DLYYC1       : in    std_ulogic;
    DLYYC2       : in    std_ulogic;
    DLYYC3       : in    std_ulogic;
    DLYYC4       : in    std_ulogic;
    DLYGLC0      : in    std_ulogic;
    DLYGLC1      : in    std_ulogic;
    DLYGLC2      : in    std_ulogic;
    DLYGLC3      : in    std_ulogic;
    DLYGLC4      : in    std_ulogic;
    FINDIV0      : in    std_ulogic;
    FINDIV1      : in    std_ulogic;
    FINDIV2      : in    std_ulogic;
    FINDIV3      : in    std_ulogic;
    FINDIV4      : in    std_ulogic;
    FINDIV5      : in    std_ulogic;
    FINDIV6      : in    std_ulogic;
    FBDIV0       : in    std_ulogic;
    FBDIV1       : in    std_ulogic;
    FBDIV2       : in    std_ulogic;
    FBDIV3       : in    std_ulogic;
    FBDIV4       : in    std_ulogic;
    FBDIV5       : in    std_ulogic;
    FBDIV6       : in    std_ulogic;
    FBDLY0       : in    std_ulogic;
    FBDlY1       : in    std_ulogic;
    FBDLY2       : in    std_ulogic;
    FBDLY3       : in    std_ulogic;
    FBDlY4       : in    std_ulogic;
    FBSEL0       : in    std_ulogic;
    FBSEL1       : in    std_ulogic;
    XDLYSEL      : in    std_ulogic;
    VCOSEL0      : in    std_ulogic;
    VCOSEL1      : in    std_ulogic;
    VCOSEL2      : in    std_ulogic;
    GLA          : out   std_ulogic;
    LOCK         : out   std_ulogic;
    GLB          : out   std_ulogic;
    YB           : out   std_ulogic;
    GLC          : out   std_ulogic;
    YC           : out   std_ulogic
   );

  attribute VITAL_LEVEL0 of PLL_V2 : entity is TRUE;
end PLL_V2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.components.all;
use igloo.PLL_TIMING_V2;

architecture VITAL_ACT of PLL_V2 is
attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal CLKA_ipd               : std_ulogic;
  signal EXTFB_ipd              : std_ulogic;
  signal POWERDOWN_ipd          : std_ulogic;
  signal OADIV0_ipd             : std_ulogic;
  signal OADIV1_ipd             : std_ulogic;
  signal OADIV2_ipd             : std_ulogic;
  signal OADIV3_ipd             : std_ulogic;
  signal OADIV4_ipd             : std_ulogic;
  signal OAMUX0_ipd             : std_ulogic;
  signal OAMUX1_ipd             : std_ulogic;
  signal OAMUX2_ipd             : std_ulogic;
  signal DLYGLA0_ipd            : std_ulogic;
  signal DLYGLA1_ipd            : std_ulogic;
  signal DLYGLA2_ipd            : std_ulogic;
  signal DLYGLA3_ipd            : std_ulogic;
  signal DLYGLA4_ipd            : std_ulogic;
  signal OBDIV0_ipd             : std_ulogic;
  signal OBDIV1_ipd             : std_ulogic;
  signal OBDIV2_ipd             : std_ulogic;
  signal OBDIV3_ipd             : std_ulogic;
  signal OBDIV4_ipd             : std_ulogic;
  signal OBMUX0_ipd             : std_ulogic;
  signal OBMUX1_ipd             : std_ulogic;
  signal OBMUX2_ipd             : std_ulogic;
  signal DLYYB0_ipd             : std_ulogic;
  signal DLYYB1_ipd             : std_ulogic;
  signal DLYYB2_ipd             : std_ulogic;
  signal DLYYB3_ipd             : std_ulogic;
  signal DLYYB4_ipd             : std_ulogic;
  signal DLYGLB0_ipd            : std_ulogic;
  signal DLYGLB1_ipd            : std_ulogic;
  signal DLYGLB2_ipd            : std_ulogic;
  signal DLYGLB3_ipd            : std_ulogic;
  signal DLYGLB4_ipd            : std_ulogic;
  signal OCDIV0_ipd             : std_ulogic;
  signal OCDIV1_ipd             : std_ulogic;
  signal OCDIV2_ipd             : std_ulogic;
  signal OCDIV3_ipd             : std_ulogic;
  signal OCDIV4_ipd             : std_ulogic;
  signal OCMUX0_ipd             : std_ulogic;
  signal OCMUX1_ipd             : std_ulogic;
  signal OCMUX2_ipd             : std_ulogic;
  signal DLYYC0_ipd             : std_ulogic;
  signal DLYYC1_ipd             : std_ulogic;
  signal DLYYC2_ipd             : std_ulogic;
  signal DLYYC3_ipd             : std_ulogic;
  signal DLYYC4_ipd             : std_ulogic;
  signal DLYGLC0_ipd            : std_ulogic;
  signal DLYGLC1_ipd            : std_ulogic;
  signal DLYGLC2_ipd            : std_ulogic;
  signal DLYGLC3_ipd            : std_ulogic;
  signal DLYGLC4_ipd            : std_ulogic;
  signal FINDIV0_ipd            : std_ulogic;
  signal FINDIV1_ipd            : std_ulogic;
  signal FINDIV2_ipd            : std_ulogic;
  signal FINDIV3_ipd            : std_ulogic;
  signal FINDIV4_ipd            : std_ulogic;
  signal FINDIV5_ipd            : std_ulogic;
  signal FINDIV6_ipd            : std_ulogic;
  signal FBDIV0_ipd             : std_ulogic;
  signal FBDIV1_ipd             : std_ulogic;
  signal FBDIV2_ipd             : std_ulogic;
  signal FBDIV3_ipd             : std_ulogic;
  signal FBDIV4_ipd             : std_ulogic;
  signal FBDIV5_ipd             : std_ulogic;
  signal FBDIV6_ipd             : std_ulogic;
  signal FBDLY0_ipd             : std_ulogic;
  signal FBDlY1_ipd             : std_ulogic;
  signal FBDLY2_ipd             : std_ulogic;
  signal FBDLY3_ipd             : std_ulogic;
  signal FBDlY4_ipd             : std_ulogic;
  signal FBSEL0_ipd             : std_ulogic;
  signal FBSEL1_ipd             : std_ulogic;
  signal XDLYSEL_ipd            : std_ulogic;
  signal VCOSEL0_ipd            : std_ulogic;
  signal VCOSEL1_ipd            : std_ulogic;
  signal VCOSEL2_ipd            : std_ulogic;

  signal GND                    : std_logic := '0';
  signal UNUSED                 : std_logic := 'X';

  component PLLPRIM
    generic (
              VCOFREQUENCY          : Real;
              f_CLKA_LOCK           : Integer;
              EMULATED_SYSTEM_DELAY : Time;
              IN_DIV_DELAY          : Time;
              OUT_DIV_DELAY         : Time;
              MUX_DELAY             : Time;
              IN_DELAY_BYP1         : Time;
              BYP_MUX_DELAY         : Time;
              GL_DRVR_DELAY         : Time;
              Y_DRVR_DELAY          : Time;
              FB_MUX_DELAY          : Time;
              X_MUX_DELAY           : Time;
              FIN_LOCK_DELAY        : Time;
              LOCK_OUT_DELAY        : Time;
              PROG_INIT_DELAY       : Time;
              PROG_STEP_INCREMENT   : Time;
              BYP0_CLK_GL           : Time;
              CLKA_TO_REF_DELAY     : Time
            );
    port (
           DYNSYNC      : in    std_ulogic;
           CLKA         : in    std_ulogic;
           EXTFB        : in    std_ulogic;
           POWERDOWN    : in    std_ulogic;
           CLKB         : in    std_ulogic;
           CLKC         : in    std_ulogic;
           OADIVRST     : in    std_ulogic;
           OADIVHALF    : in    std_ulogic;
           OADIV0       : in    std_ulogic;
           OADIV1       : in    std_ulogic;
           OADIV2       : in    std_ulogic;
           OADIV3       : in    std_ulogic;
           OADIV4       : in    std_ulogic;
           OAMUX0       : in    std_ulogic;
           OAMUX1       : in    std_ulogic;
           OAMUX2       : in    std_ulogic;
           DLYGLA0      : in    std_ulogic;
           DLYGLA1      : in    std_ulogic;
           DLYGLA2      : in    std_ulogic;
           DLYGLA3      : in    std_ulogic;
           DLYGLA4      : in    std_ulogic;
           OBDIVRST     : in    std_ulogic;
           OBDIVHALF    : in    std_ulogic;
           OBDIV0       : in    std_ulogic;
           OBDIV1       : in    std_ulogic;
           OBDIV2       : in    std_ulogic;
           OBDIV3       : in    std_ulogic;
           OBDIV4       : in    std_ulogic;
           OBMUX0       : in    std_ulogic;
           OBMUX1       : in    std_ulogic;
           OBMUX2       : in    std_ulogic;
           DLYYB0       : in    std_ulogic;
           DLYYB1       : in    std_ulogic;
           DLYYB2       : in    std_ulogic;
           DLYYB3       : in    std_ulogic;
           DLYYB4       : in    std_ulogic;
           DLYGLB0      : in    std_ulogic;
           DLYGLB1      : in    std_ulogic;
           DLYGLB2      : in    std_ulogic;
           DLYGLB3      : in    std_ulogic;
           DLYGLB4      : in    std_ulogic;
           OCDIVRST     : in    std_ulogic;
           OCDIVHALF    : in    std_ulogic;
           OCDIV0       : in    std_ulogic;
           OCDIV1       : in    std_ulogic;
           OCDIV2       : in    std_ulogic;
           OCDIV3       : in    std_ulogic;
           OCDIV4       : in    std_ulogic;
           OCMUX0       : in    std_ulogic;
           OCMUX1       : in    std_ulogic;
           OCMUX2       : in    std_ulogic;
           DLYYC0       : in    std_ulogic;
           DLYYC1       : in    std_ulogic;
           DLYYC2       : in    std_ulogic;
           DLYYC3       : in    std_ulogic;
           DLYYC4       : in    std_ulogic;
           DLYGLC0      : in    std_ulogic;
           DLYGLC1      : in    std_ulogic;
           DLYGLC2      : in    std_ulogic;
           DLYGLC3      : in    std_ulogic;
           DLYGLC4      : in    std_ulogic;
           FINDIV0      : in    std_ulogic;
           FINDIV1      : in    std_ulogic;
           FINDIV2      : in    std_ulogic;
           FINDIV3      : in    std_ulogic;
           FINDIV4      : in    std_ulogic;
           FINDIV5      : in    std_ulogic;
           FINDIV6      : in    std_ulogic;
           FBDIV0       : in    std_ulogic;
           FBDIV1       : in    std_ulogic;
           FBDIV2       : in    std_ulogic;
           FBDIV3       : in    std_ulogic;
           FBDIV4       : in    std_ulogic;
           FBDIV5       : in    std_ulogic;
           FBDIV6       : in    std_ulogic;
           FBDLY0       : in    std_ulogic;
           FBDlY1       : in    std_ulogic;
           FBDLY2       : in    std_ulogic;
           FBDLY3       : in    std_ulogic;
           FBDlY4       : in    std_ulogic;
           FBSEL0       : in    std_ulogic;
           FBSEL1       : in    std_ulogic;
           XDLYSEL      : in    std_ulogic;
           VCOSEL0      : in    std_ulogic;
           VCOSEL1      : in    std_ulogic;
           VCOSEL2      : in    std_ulogic;
           GLA          : out   std_ulogic;
           LOCK         : out   std_ulogic;
           GLB          : out   std_ulogic;
           YB           : out   std_ulogic;
           GLC          : out   std_ulogic;
           YC           : out   std_ulogic
         );
  end component;

  begin

    ---------------------
    --  INPUT PATH DELAYs
    ---------------------
    WireDelay : block

    begin

      VitalWireDelay ( CLKA_ipd,      CLKA,      tipd_CLKA );
      VitalWireDelay ( EXTFB_ipd,     EXTFB,     tipd_EXTFB );
      VitalWireDelay ( POWERDOWN_ipd, POWERDOWN, tipd_POWERDOWN );
      VitalWireDelay ( OADIV0_ipd,    OADIV0,    tipd_OADIV0 );
      VitalWireDelay ( OADIV1_ipd,    OADIV1,    tipd_OADIV1 );
      VitalWireDelay ( OADIV2_ipd,    OADIV2,    tipd_OADIV2 );
      VitalWireDelay ( OADIV3_ipd,    OADIV3,    tipd_OADIV3 );
      VitalWireDelay ( OADIV4_ipd,    OADIV4,    tipd_OADIV4 );
      VitalWireDelay ( OAMUX0_ipd,    OAMUX0,    tipd_OAMUX0 );
      VitalWireDelay ( OAMUX1_ipd,    OAMUX1,    tipd_OAMUX1 );
      VitalWireDelay ( OAMUX2_ipd,    OAMUX2,    tipd_OAMUX2 );
      VitalWireDelay ( DLYGLA0_ipd,   DLYGLA0,   tipd_DLYGLA0 );
      VitalWireDelay ( DLYGLA1_ipd,   DLYGLA1,   tipd_DLYGLA1 );
      VitalWireDelay ( DLYGLA2_ipd,   DLYGLA2,   tipd_DLYGLA2 );
      VitalWireDelay ( DLYGLA3_ipd,   DLYGLA3,   tipd_DLYGLA3 );
      VitalWireDelay ( DLYGLA4_ipd,   DLYGLA4,   tipd_DLYGLA4 );
      VitalWireDelay ( OBDIV0_ipd,    OBDIV0,    tipd_OBDIV0 );
      VitalWireDelay ( OBDIV1_ipd,    OBDIV1,    tipd_OBDIV1 );
      VitalWireDelay ( OBDIV2_ipd,    OBDIV2,    tipd_OBDIV2 );
      VitalWireDelay ( OBDIV3_ipd,    OBDIV3,    tipd_OBDIV3 );
      VitalWireDelay ( OBDIV4_ipd,    OBDIV4,    tipd_OBDIV4 );
      VitalWireDelay ( OBMUX0_ipd,    OBMUX0,    tipd_OBMUX0 );
      VitalWireDelay ( OBMUX1_ipd,    OBMUX1,    tipd_OBMUX1 );
      VitalWireDelay ( OBMUX2_ipd,    OBMUX2,    tipd_OBMUX2 );
      VitalWireDelay ( DLYYB0_ipd,    DLYYB0,    tipd_DLYYB0 );
      VitalWireDelay ( DLYYB1_ipd,    DLYYB1,    tipd_DLYYB1 );
      VitalWireDelay ( DLYYB2_ipd,    DLYYB2,    tipd_DLYYB2 );
      VitalWireDelay ( DLYYB3_ipd,    DLYYB3,    tipd_DLYYB3 );
      VitalWireDelay ( DLYYB4_ipd,    DLYYB4,    tipd_DLYYB4 );
      VitalWireDelay ( DLYGLB0_ipd,   DLYGLB0,   tipd_DLYGLB0 );
      VitalWireDelay ( DLYGLB1_ipd,   DLYGLB1,   tipd_DLYGLB1 );
      VitalWireDelay ( DLYGLB2_ipd,   DLYGLB2,   tipd_DLYGLB2 );
      VitalWireDelay ( DLYGLB3_ipd,   DLYGLB3,   tipd_DLYGLB3 );
      VitalWireDelay ( DLYGLB4_ipd,   DLYGLB4,   tipd_DLYGLB4 );
      VitalWireDelay ( OCDIV0_ipd,    OCDIV0,    tipd_OCDIV0 );
      VitalWireDelay ( OCDIV1_ipd,    OCDIV1,    tipd_OCDIV1 );
      VitalWireDelay ( OCDIV2_ipd,    OCDIV2,    tipd_OCDIV2 );
      VitalWireDelay ( OCDIV3_ipd,    OCDIV3,    tipd_OCDIV3 );
      VitalWireDelay ( OCDIV4_ipd,    OCDIV4,    tipd_OCDIV4 );
      VitalWireDelay ( OCMUX0_ipd,    OCMUX0,    tipd_OCMUX0 );
      VitalWireDelay ( OCMUX1_ipd,    OCMUX1,    tipd_OCMUX1 );
      VitalWireDelay ( OCMUX2_ipd,    OCMUX2,    tipd_OCMUX2 );
      VitalWireDelay ( DLYYC0_ipd,    DLYYC0,    tipd_DLYYC0 );
      VitalWireDelay ( DLYYC1_ipd,    DLYYC1,    tipd_DLYYC1 );
      VitalWireDelay ( DLYYC2_ipd,    DLYYC2,    tipd_DLYYC2 );
      VitalWireDelay ( DLYYC3_ipd,    DLYYC3,    tipd_DLYYC3 );
      VitalWireDelay ( DLYYC4_ipd,    DLYYC4,    tipd_DLYYC4 );
      VitalWireDelay ( DLYGLC0_ipd,   DLYGLC0,   tipd_DLYGLC0 );
      VitalWireDelay ( DLYGLC1_ipd,   DLYGLC1,   tipd_DLYGLC1 );
      VitalWireDelay ( DLYGLC2_ipd,   DLYGLC2,   tipd_DLYGLC2 );
      VitalWireDelay ( DLYGLC3_ipd,   DLYGLC3,   tipd_DLYGLC3 );
      VitalWireDelay ( DLYGLC4_ipd,   DLYGLC4,   tipd_DLYGLC4 );
      VitalWireDelay ( FINDIV0_ipd,   FINDIV0,   tipd_FINDIV0 );
      VitalWireDelay ( FINDIV1_ipd,   FINDIV1,   tipd_FINDIV1 );
      VitalWireDelay ( FINDIV2_ipd,   FINDIV2,   tipd_FINDIV2 );
      VitalWireDelay ( FINDIV3_ipd,   FINDIV3,   tipd_FINDIV3 );
      VitalWireDelay ( FINDIV4_ipd,   FINDIV4,   tipd_FINDIV4 );
      VitalWireDelay ( FINDIV5_ipd,   FINDIV5,   tipd_FINDIV5 );
      VitalWireDelay ( FINDIV6_ipd,   FINDIV6,   tipd_FINDIV6 );
      VitalWireDelay ( FBDIV0_ipd,    FBDIV0,    tipd_FBDIV0 );
      VitalWireDelay ( FBDIV1_ipd,    FBDIV1,    tipd_FBDIV1 );
      VitalWireDelay ( FBDIV2_ipd,    FBDIV2,    tipd_FBDIV2 );
      VitalWireDelay ( FBDIV3_ipd,    FBDIV3,    tipd_FBDIV3 );
      VitalWireDelay ( FBDIV4_ipd,    FBDIV4,    tipd_FBDIV4 );
      VitalWireDelay ( FBDIV5_ipd,    FBDIV5,    tipd_FBDIV5 );
      VitalWireDelay ( FBDIV6_ipd,    FBDIV6,    tipd_FBDIV6 );
      VitalWireDelay ( FBDLY0_ipd,    FBDLY0,    tipd_FBDLY0 );
      VitalWireDelay ( FBDLY1_ipd,    FBDLY1,    tipd_FBDLY1 );
      VitalWireDelay ( FBDLY2_ipd,    FBDLY2,    tipd_FBDLY2 );
      VitalWireDelay ( FBDLY3_ipd,    FBDLY3,    tipd_FBDLY3 );
      VitalWireDelay ( FBDLY4_ipd,    FBDLY4,    tipd_FBDLY4 );
      VitalWireDelay ( FBSEL0_ipd,    FBSEL0,    tipd_FBSEL0 );
      VitalWireDelay ( FBSEL1_ipd,    FBSEL1,    tipd_FBSEL1 );
      VitalWireDelay ( XDLYSEL_ipd,   XDLYSEL,   tipd_XDLYSEL );
      VitalWireDelay ( VCOSEL0_ipd,   VCOSEL0,   tipd_VCOSEL0 );
      VitalWireDelay ( VCOSEL1_ipd,   VCOSEL1,   tipd_VCOSEL1 );
      VitalWireDelay ( VCOSEL2_ipd,   VCOSEL2,   tipd_VCOSEL2 );
 
    end block WireDelay;
    
    P1: PLLPRIM
          generic map (
                        VCOFREQUENCY          => VCOFREQUENCY,
                        f_CLKA_LOCK           => f_CLKA_LOCK,
                        EMULATED_SYSTEM_DELAY => PLL_TIMING_V2.EMULATED_SYSTEM_DELAY,
                        IN_DIV_DELAY          => PLL_TIMING_V2.IN_DIV_DELAY,
                        OUT_DIV_DELAY         => PLL_TIMING_V2.OUT_DIV_DELAY,
                        MUX_DELAY             => PLL_TIMING_V2.MUX_DELAY,
                        IN_DELAY_BYP1         => PLL_TIMING_V2.IN_DELAY_BYP1,
                        BYP_MUX_DELAY         => PLL_TIMING_V2.BYP_MUX_DELAY,
                        GL_DRVR_DELAY         => PLL_TIMING_V2.GL_DRVR_DELAY,
                        Y_DRVR_DELAY          => PLL_TIMING_V2.Y_DRVR_DELAY,
                        FB_MUX_DELAY          => PLL_TIMING_V2.FB_MUX_DELAY,
                        X_MUX_DELAY           => PLL_TIMING_V2.X_MUX_DELAY,
                        FIN_LOCK_DELAY        => PLL_TIMING_V2.FIN_LOCK_DELAY,
                        LOCK_OUT_DELAY        => PLL_TIMING_V2.LOCK_OUT_DELAY,
                        PROG_INIT_DELAY       => PLL_TIMING_V2.PROG_INIT_DELAY,
                        PROG_STEP_INCREMENT   => PLL_TIMING_V2.PROG_STEP_INCREMENT,
                        BYP0_CLK_GL           => PLL_TIMING_V2.BYP0_CLK_GL,
                        CLKA_TO_REF_DELAY     => PLL_TIMING_V2.CLKA_TO_REF_DELAY
                      )
          port map    (
                        DYNSYNC      => GND,
                        CLKA         => CLKA_ipd,
                        EXTFB        => EXTFB_ipd,
                        POWERDOWN    => POWERDOWN_ipd,
                        CLKB         => UNUSED,
                        CLKC         => UNUSED,
                        OADIVRST     => GND,
                        OADIVHALF    => GND,
                        OADIV0       => OADIV0_ipd,
                        OADIV1       => OADIV1_ipd,
                        OADIV2       => OADIV2_ipd,
                        OADIV3       => OADIV3_ipd,
                        OADIV4       => OADIV4_ipd,
                        OAMUX0       => OAMUX0_ipd,
                        OAMUX1       => OAMUX1_ipd,
                        OAMUX2       => OAMUX2_ipd,
                        DLYGLA0      => DLYGLA0_ipd,
                        DLYGLA1      => DLYGLA1_ipd,
                        DLYGLA2      => DLYGLA2_ipd,
                        DLYGLA3      => DLYGLA3_ipd,
                        DLYGLA4      => DLYGLA4_ipd,
                        OBDIVRST     => GND,
                        OBDIVHALF    => GND,
                        OBDIV0       => OBDIV0_ipd,
                        OBDIV1       => OBDIV1_ipd,
                        OBDIV2       => OBDIV2_ipd,
                        OBDIV3       => OBDIV3_ipd,
                        OBDIV4       => OBDIV4_ipd,
                        OBMUX0       => OBMUX0_ipd,
                        OBMUX1       => OBMUX1_ipd,
                        OBMUX2       => OBMUX2_ipd,
                        DLYYB0       => DLYYB0_ipd,
                        DLYYB1       => DLYYB1_ipd,
                        DLYYB2       => DLYYB2_ipd,
                        DLYYB3       => DLYYB3_ipd,
                        DLYYB4       => DLYYB4_ipd,
                        DLYGLB0      => DLYGLB0_ipd,
                        DLYGLB1      => DLYGLB1_ipd,
                        DLYGLB2      => DLYGLB2_ipd,
                        DLYGLB3      => DLYGLB3_ipd,
                        DLYGLB4      => DLYGLB4_ipd,
                        OCDIVRST     => GND,
                        OCDIVHALF    => GND,
                        OCDIV0       => OCDIV0_ipd,
                        OCDIV1       => OCDIV1_ipd,
                        OCDIV2       => OCDIV2_ipd,
                        OCDIV3       => OCDIV3_ipd,
                        OCDIV4       => OCDIV4_ipd,
                        OCMUX0       => OCMUX0_ipd,
                        OCMUX1       => OCMUX1_ipd,
                        OCMUX2       => OCMUX2_ipd,
                        DLYYC0       => DLYYC0_ipd,
                        DLYYC1       => DLYYC1_ipd,
                        DLYYC2       => DLYYC2_ipd,
                        DLYYC3       => DLYYC3_ipd,
                        DLYYC4       => DLYYC4_ipd,
                        DLYGLC0      => DLYGLC0_ipd,
                        DLYGLC1      => DLYGLC1_ipd,
                        DLYGLC2      => DLYGLC2_ipd,
                        DLYGLC3      => DLYGLC3_ipd,
                        DLYGLC4      => DLYGLC4_ipd,
                        FINDIV0      => FINDIV0_ipd,
                        FINDIV1      => FINDIV1_ipd,
                        FINDIV2      => FINDIV2_ipd,
                        FINDIV3      => FINDIV3_ipd,
                        FINDIV4      => FINDIV4_ipd,
                        FINDIV5      => FINDIV5_ipd,
                        FINDIV6      => FINDIV6_ipd,
                        FBDIV0       => FBDIV0_ipd,
                        FBDIV1       => FBDIV1_ipd,
                        FBDIV2       => FBDIV2_ipd,
                        FBDIV3       => FBDIV3_ipd,
                        FBDIV4       => FBDIV4_ipd,
                        FBDIV5       => FBDIV5_ipd,
                        FBDIV6       => FBDIV6_ipd,
                        FBDLY0       => FBDLY0_ipd,
                        FBDlY1       => FBDlY1_ipd,
                        FBDLY2       => FBDLY2_ipd,
                        FBDLY3       => FBDLY3_ipd,
                        FBDlY4       => FBDlY4_ipd,
                        FBSEL0       => FBSEL0_ipd,
                        FBSEL1       => FBSEL1_ipd,
                        XDLYSEL      => XDLYSEL_ipd,
                        VCOSEL0      => VCOSEL0_ipd,
                        VCOSEL1      => VCOSEL1_ipd,
                        VCOSEL2      => VCOSEL2_ipd,
                        GLA          => GLA,
                        LOCK         => LOCK,
                        GLB          => GLB,
                        YB           => YB,
                        GLC          => GLC,
                        YC           => YC
                      );

  end VITAL_ACT;

configuration CFG_PLL_V2_VITAL of PLL_V2 is
  for VITAL_ACT
  end for;
end CFG_PLL_V2_VITAL;

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
 entity SHREG is
   generic(
      tipd_SDIN      : VitalDelayType01 := ( 0.0 ns, 0.0 ns );
      tipd_SCLK      : VitalDelayType01 := ( 0.0 ns, 0.0 ns );
      tipd_SSHIFT    : VitalDelayType01 := ( 0.0 ns, 0.0 ns );
      tipd_SUPDATE   : VitalDelayType01 := ( 0.0 ns, 0.0 ns );

      TimingChecksOn : Boolean := True;
      InstancePath   : STRING  := "*";
      Xon            : Boolean := False;
      MsgOn          : Boolean := True);

   port(
      SDIN           :	in    STD_ULOGIC; -- Serial data input
      SCLK           :	in    STD_ULOGIC; -- Serial Clock signal
      SSHIFT         :	in    STD_ULOGIC; -- Serial shift enable signal 
      SUPDATE        :	in    STD_ULOGIC; -- Data in SR loaded into update latch
      SDOUT          :	out   STD_ULOGIC; -- Serial data output - data from LSB of SR shifted out
      SUPDATELATCH   :  out   STD_LOGIC_VECTOR ( 80 downto 0 )); -- Configuration bits

attribute VITAL_LEVEL0 of SHREG : entity is TRUE;
end SHREG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of SHREG is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL SDIN_ipd    : STD_ULOGIC := 'X';
   SIGNAL SCLK_ipd    : STD_ULOGIC := 'X';
   SIGNAL SSHIFT_ipd  : STD_ULOGIC := 'X';
   SIGNAL SUPDATE_ipd : STD_ULOGIC := 'X';

   SIGNAL SH_REG      : STD_LOGIC_VECTOR ( 80 downto 0 ) := ( OTHERS => 'X' );

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

     VitalWireDelay ( SDIN_ipd,    SDIN,    tipd_SDIN );
     VitalWireDelay ( SCLK_ipd,    SCLK,    tipd_SCLK );
     VitalWireDelay ( SSHIFT_ipd,  SSHIFT,  tipd_SSHIFT );
     VitalWireDelay ( SUPDATE_ipd, SUPDATE, tipd_SUPDATE );

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process ( SCLK_ipd )

  begin

    if ( SCLK_ipd'event and ( TO_X01 ( SCLK_ipd ) = '1' )) then
      if ( TO_X01 ( SSHIFT_ipd ) = '1' ) then
        SH_REG <= SDIN_ipd & SH_REG ( 80 downto 1 );
        SDOUT <= SH_REG ( 0 );
      else
        SH_REG <= SH_REG ( 80 downto 0 );
      end if;
    end if;

  end process VITALBehavior;

  VITALBehavior2: process ( SUPDATE_ipd, SH_REG )
  begin
    if ( TO_X01 ( SUPDATE_ipd ) = '1' ) then   
       SUPDATELATCH <= SH_REG ( 80 downto 0 );
    end if;
  end process VITALBehavior2;


end VITAL_ACT;

configuration CFG_SHREG_VITAL of SHREG is
  for VITAL_ACT
  end for;
end CFG_SHREG_VITAL;

library IEEE;
use IEEE.VITAL_Timing.all;
use IEEE.STD_LOGIC_1164.all;

-- SHREG shifts in 81 bits, but only bits 79 - 0 are included in the  
-- configuration bit string.  Bit 80 used as the RESET ENABLE.  Bits
-- 71 - 73 and 77 - 49 not used by simulation model.

-- entity declaration --
 entity DYNCCC is
   generic(
      VCOFREQUENCY      :  Real    := 0.0;
      f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

      TimingChecksOn    :  Boolean := True;
      InstancePath      :  STRING  := "*";
      Xon               :  Boolean := False;
      MsgOn             :  Boolean := True;

      tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKC         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SDIN         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SCLK         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SSHIFT       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SUPDATE      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_MODE         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

      tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );

      tpd_SCLK_SDOUT    : VitalDelayType01  := ( 0.100 ns, 0.100 ns );

      tsetup_SSHIFT_SCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_SSHIFT_SCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_negedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_SDIN_SCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_SDIN_SCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_negedge_posedge    : VitalDelayType := 0.000 ns;

      tpw_SUPDATE_posedge                : VitalDelayType := 0.000 ns; 
      tpw_SUPDATE_negedge                : VitalDelayType := 0.000 ns; 
      tpw_SCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_SCLK_negedge                   : VitalDelayType := 0.000 ns

      ); 

   port (
          CLKA         : in    std_ulogic;
          EXTFB        : in    std_ulogic;
          POWERDOWN    : in    std_ulogic;
          CLKB         : in    std_ulogic;
          CLKC         : in    std_ulogic;
          SDIN         : in    std_ulogic;
          SCLK         : in    std_ulogic;
          SSHIFT       : in    std_ulogic;
          SUPDATE      : in    std_ulogic;
          MODE         : in    std_ulogic;
          OADIV0       : in    std_ulogic;
          OADIV1       : in    std_ulogic;
          OADIV2       : in    std_ulogic;
          OADIV3       : in    std_ulogic;
          OADIV4       : in    std_ulogic;
          OAMUX0       : in    std_ulogic;
          OAMUX1       : in    std_ulogic;
          OAMUX2       : in    std_ulogic;
          DLYGLA0      : in    std_ulogic;
          DLYGLA1      : in    std_ulogic;
          DLYGLA2      : in    std_ulogic;
          DLYGLA3      : in    std_ulogic;
          DLYGLA4      : in    std_ulogic;
          OBDIV0       : in    std_ulogic;
          OBDIV1       : in    std_ulogic;
          OBDIV2       : in    std_ulogic;
          OBDIV3       : in    std_ulogic;
          OBDIV4       : in    std_ulogic;
          OBMUX0       : in    std_ulogic;
          OBMUX1       : in    std_ulogic;
          OBMUX2       : in    std_ulogic;
          DLYYB0       : in    std_ulogic;
          DLYYB1       : in    std_ulogic;
          DLYYB2       : in    std_ulogic;
          DLYYB3       : in    std_ulogic;
          DLYYB4       : in    std_ulogic;
          DLYGLB0      : in    std_ulogic;
          DLYGLB1      : in    std_ulogic;
          DLYGLB2      : in    std_ulogic;
          DLYGLB3      : in    std_ulogic;
          DLYGLB4      : in    std_ulogic;
          OCDIV0       : in    std_ulogic;
          OCDIV1       : in    std_ulogic;
          OCDIV2       : in    std_ulogic;
          OCDIV3       : in    std_ulogic;
          OCDIV4       : in    std_ulogic;
          OCMUX0       : in    std_ulogic;
          OCMUX1       : in    std_ulogic;
          OCMUX2       : in    std_ulogic;
          DLYYC0       : in    std_ulogic;
          DLYYC1       : in    std_ulogic;
          DLYYC2       : in    std_ulogic;
          DLYYC3       : in    std_ulogic;
          DLYYC4       : in    std_ulogic;
          DLYGLC0      : in    std_ulogic;
          DLYGLC1      : in    std_ulogic;
          DLYGLC2      : in    std_ulogic;
          DLYGLC3      : in    std_ulogic;
          DLYGLC4      : in    std_ulogic;
          FINDIV0      : in    std_ulogic;
          FINDIV1      : in    std_ulogic;
          FINDIV2      : in    std_ulogic;
          FINDIV3      : in    std_ulogic;
          FINDIV4      : in    std_ulogic;
          FINDIV5      : in    std_ulogic;
          FINDIV6      : in    std_ulogic;
          FBDIV0       : in    std_ulogic;
          FBDIV1       : in    std_ulogic;
          FBDIV2       : in    std_ulogic;
          FBDIV3       : in    std_ulogic;
          FBDIV4       : in    std_ulogic;
          FBDIV5       : in    std_ulogic;
          FBDIV6       : in    std_ulogic;
          FBDLY0       : in    std_ulogic;
          FBDlY1       : in    std_ulogic;
          FBDLY2       : in    std_ulogic;
          FBDLY3       : in    std_ulogic;
          FBDlY4       : in    std_ulogic;
          FBSEL0       : in    std_ulogic;
          FBSEL1       : in    std_ulogic;
          XDLYSEL      : in    std_ulogic;
          VCOSEL0      : in    std_ulogic;
          VCOSEL1      : in    std_ulogic;
          VCOSEL2      : in    std_ulogic;
          GLA          : out   std_ulogic;
          LOCK         : out   std_ulogic;
          GLB          : out   std_ulogic;
          YB           : out   std_ulogic;
          GLC          : out   std_ulogic;
          YC           : out   std_ulogic;
          SDOUT        : out   std_ulogic
        );

attribute VITAL_LEVEL0 of DYNCCC : entity is TRUE;
end DYNCCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.components.all;

architecture VITAL_ACT of DYNCCC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal CLKA_ipd               : std_ulogic;
   signal EXTFB_ipd              : std_ulogic;
   signal POWERDOWN_ipd          : std_ulogic;
   signal CLKB_ipd               : std_ulogic;
   signal CLKC_ipd               : std_ulogic;
   signal SDIN_ipd               : std_ulogic;
   signal SCLK_ipd               : std_ulogic;
   signal SSHIFT_ipd             : std_ulogic;
   signal SUPDATE_ipd            : std_ulogic;
   signal MODE_ipd               : std_ulogic;

   signal C            : std_logic_vector ( 79 downto 0 ) := ( others => 'X' );
   signal SUPDATELATCH : std_logic_vector ( 80 downto 0 ) := ( others => 'X' );
   signal PC           : std_logic_vector ( 79 downto 0 ) := ( others => 'X' );

   -- Unused configuration bits
   signal DYNCSEL                : std_ulogic;
   signal DYNBSEL                : std_ulogic;
   signal DYNASEL                : std_ulogic;
   signal STATCSEL               : std_ulogic;
   signal STATBSEL               : std_ulogic;
   signal STATASEL               : std_ulogic;

   -- SDOUT SHREG port map
   signal SDOUT_zd               : std_ulogic;

   -- synchronisation trigger generated based on SUPDATE, MODE and SUPDATELATCH(80)
   signal DYNSYNC                : std_ulogic := '0';

   signal GND                    : std_logic  := '0';

   component PLLPRIM
     generic (
              VCOFREQUENCY :  Real;
              f_CLKA_LOCK  :  Integer
             );
     port (
            DYNSYNC      : in    std_ulogic;
            CLKA         : in    std_ulogic;
            EXTFB        : in    std_ulogic;
            POWERDOWN    : in    std_ulogic;
            CLKB         : in    std_ulogic;
            CLKC         : in    std_ulogic;
            OADIVRST     : in    std_ulogic;
            OADIVHALF    : in    std_ulogic;
            OADIV0       : in    std_ulogic;
            OADIV1       : in    std_ulogic;
            OADIV2       : in    std_ulogic;
            OADIV3       : in    std_ulogic;
            OADIV4       : in    std_ulogic;
            OAMUX0       : in    std_ulogic;
            OAMUX1       : in    std_ulogic;
            OAMUX2       : in    std_ulogic;
            DLYGLA0      : in    std_ulogic;
            DLYGLA1      : in    std_ulogic;
            DLYGLA2      : in    std_ulogic;
            DLYGLA3      : in    std_ulogic;
            DLYGLA4      : in    std_ulogic;
            OBDIVRST     : in    std_ulogic;
            OBDIVHALF    : in    std_ulogic;
            OBDIV0       : in    std_ulogic;
            OBDIV1       : in    std_ulogic;
            OBDIV2       : in    std_ulogic;
            OBDIV3       : in    std_ulogic;
            OBDIV4       : in    std_ulogic;
            OBMUX0       : in    std_ulogic;
            OBMUX1       : in    std_ulogic;
            OBMUX2       : in    std_ulogic;
            DLYYB0       : in    std_ulogic;
            DLYYB1       : in    std_ulogic;
            DLYYB2       : in    std_ulogic;
            DLYYB3       : in    std_ulogic;
            DLYYB4       : in    std_ulogic;
            DLYGLB0      : in    std_ulogic;
            DLYGLB1      : in    std_ulogic;
            DLYGLB2      : in    std_ulogic;
            DLYGLB3      : in    std_ulogic;
            DLYGLB4      : in    std_ulogic;
            OCDIVRST     : in    std_ulogic;
            OCDIVHALF    : in    std_ulogic;
            OCDIV0       : in    std_ulogic;
            OCDIV1       : in    std_ulogic;
            OCDIV2       : in    std_ulogic;
            OCDIV3       : in    std_ulogic;
            OCDIV4       : in    std_ulogic;
            OCMUX0       : in    std_ulogic;
            OCMUX1       : in    std_ulogic;
            OCMUX2       : in    std_ulogic;
            DLYYC0       : in    std_ulogic;
            DLYYC1       : in    std_ulogic;
            DLYYC2       : in    std_ulogic;
            DLYYC3       : in    std_ulogic;
            DLYYC4       : in    std_ulogic;
            DLYGLC0      : in    std_ulogic;
            DLYGLC1      : in    std_ulogic;
            DLYGLC2      : in    std_ulogic;
            DLYGLC3      : in    std_ulogic;
            DLYGLC4      : in    std_ulogic;
            FINDIV0      : in    std_ulogic;
            FINDIV1      : in    std_ulogic;
            FINDIV2      : in    std_ulogic;
            FINDIV3      : in    std_ulogic;
            FINDIV4      : in    std_ulogic;
            FINDIV5      : in    std_ulogic;
            FINDIV6      : in    std_ulogic;
            FBDIV0       : in    std_ulogic;
            FBDIV1       : in    std_ulogic;
            FBDIV2       : in    std_ulogic;
            FBDIV3       : in    std_ulogic;
            FBDIV4       : in    std_ulogic;
            FBDIV5       : in    std_ulogic;
            FBDIV6       : in    std_ulogic;
            FBDLY0       : in    std_ulogic;
            FBDlY1       : in    std_ulogic;
            FBDLY2       : in    std_ulogic;
            FBDLY3       : in    std_ulogic;
            FBDlY4       : in    std_ulogic;
            FBSEL0       : in    std_ulogic;
            FBSEL1       : in    std_ulogic;
            XDLYSEL      : in    std_ulogic;
            VCOSEL0      : in    std_ulogic;
            VCOSEL1      : in    std_ulogic;
            VCOSEL2      : in    std_ulogic;
            GLA          : out   std_ulogic;
            LOCK         : out   std_ulogic;
            GLB          : out   std_ulogic;
            YB           : out   std_ulogic;
            GLC          : out   std_ulogic;
            YC           : out   std_ulogic
          );
     end component;

     component SHREG
       port (
              SDIN           :	in    std_ulogic;
              SCLK           :	in    std_ulogic;
              SSHIFT         :	in    std_ulogic;
              SUPDATE        :	in    std_ulogic;
              SDOUT          :	out   std_ulogic;
              SUPDATELATCH   :  out   std_logic_vector ( 80 downto 0 )
            );
     end component;
    
begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

      VitalWireDelay ( CLKA_ipd,      CLKA,      tipd_CLKA      );
      VitalWireDelay ( EXTFB_ipd,     EXTFB,     tipd_EXTFB     );
      VitalWireDelay ( POWERDOWN_ipd, POWERDOWN, tipd_POWERDOWN );
      VitalWireDelay ( CLKB_ipd,      CLKB,      tipd_CLKB      );
      VitalWireDelay ( CLKC_ipd,      CLKC,      tipd_CLKC      );
      VitalWireDelay ( SDIN_ipd,      SDIN,      tipd_SDIN      );
      VitalWireDelay ( SCLK_ipd,      SCLK,      tipd_SCLK      );
      VitalWireDelay ( SSHIFT_ipd,    SSHIFT,    tipd_SSHIFT    );
      VitalWireDelay ( SUPDATE_ipd,   SUPDATE,   tipd_SUPDATE   );
      VitalWireDelay ( MODE_ipd,      MODE,      tipd_MODE      );

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  
  PC <= 
        DYNCSEL  &
        DYNBSEL  &
        DYNASEL  &
        VCOSEL2  & 
        VCOSEL1  & 
        VCOSEL0  & 
        STATCSEL &
        STATBSEL &
        STATASEL &
        DLYYC4   &
        DLYYC3   &
        DLYYC2   &
        DLYYC1   &
        DLYYC0   &
        DLYYB4   &
        DLYYB3   &
        DLYYB2   &
        DLYYB1   &
        DLYYB0   &
        DLYGLC4  &
        DLYGLC3  &
        DLYGLC2  &
        DLYGLC1  &
        DLYGLC0  &
        DLYGLB4  &
        DLYGLB3  &
        DLYGLB2  &
        DLYGLB1  &
        DLYGLB0  &
        DLYGLA4  &
        DLYGLA3  &
        DLYGLA2  &
        DLYGLA1  &
        DLYGLA0  &
        XDLYSEL  &
        FBDLY4   &
        FBDLY3   &
        FBDLY2   &
        FBDLY1   &
        FBDLY0   &
        FBSEL1   &
        FBSEL0   &
        OCMUX2   &
        OCMUX1   &
        OCMUX0   &
        OBMUX2   &
        OBMUX1   &
        OBMUX0   &
        OAMUX2   &
        OAMUX1   &
        OAMUX0   &
        OCDIV4   &
        OCDIV3   &
        OCDIV2   &
        OCDIV1   &
        OCDIV0   &
        OBDIV4   &
        OBDIV3   &
        OBDIV2   &
        OBDIV1   &
        OBDIV0   &
        OADIV4   &
        OADIV3   &
        OADIV2   &
        OADIV1   &
        OADIV0   &
        FBDIV6   &
        FBDIV5   &
        FBDIV4   &
        FBDIV3   &
        FBDIV2   &
        FBDIV1   &
        FBDIV0   &
        FINDIV6  &
        FINDIV5  &
        FINDIV4  &
        FINDIV3  &
        FINDIV2  &
        FINDIV1  &
        FINDIV0  ;

  C <= SUPDATELATCH ( 79 downto 0 ) when ( TO_X01 ( MODE_ipd ) = '1' ) else
       PC ( 79 downto 0 ) when ( TO_X01 ( MODE_ipd ) = '0' ) else
       "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";

  -- logic for generating DYNSYNC

  latch_mode_reset : process ( SUPDATE_ipd )

    variable RESETENA_latched : std_ulogic;

  begin

    if ( TO_X01 ( SUPDATE_ipd ) = '1' ) then
      if ( TO_X01( MODE_ipd ) = '1' and TO_X01( RESETENA_latched ) = '1' ) then
        DYNSYNC <= '1'; 
      end if;
    elsif ( TO_X01 ( SUPDATE_ipd ) = '0' ) then
      DYNSYNC <= '0';
      RESETENA_latched := SUPDATELATCH ( 80 );
    end if;

  end process;


  P1: PLLPRIM 
      generic map (
                    VCOFREQUENCY => VCOFREQUENCY,
                    f_CLKA_LOCK  => f_CLKA_LOCK
                  )
      port map    ( 
                    DYNSYNC      => DYNSYNC,
                    CLKA         => CLKA_ipd,
                    EXTFB        => EXTFB_ipd,
                    POWERDOWN    => POWERDOWN_ipd,
                    CLKB         => CLKB_ipd,
                    CLKC         => CLKC_ipd,
                    OADIVRST     => GND,
                    OADIVHALF    => GND,
                    OADIV0       => C ( 14 ),
                    OADIV1       => C ( 15 ),
                    OADIV2       => C ( 16 ),
                    OADIV3       => C ( 17 ),
                    OADIV4       => C ( 18 ),
                    OAMUX0       => C ( 29 ),
                    OAMUX1       => C ( 30 ),
                    OAMUX2       => C ( 31 ),
                    DLYGLA0      => C ( 46 ),
                    DLYGLA1      => C ( 47 ),
                    DLYGLA2      => C ( 48 ),
                    DLYGLA3      => C ( 49 ),
                    DLYGLA4      => C ( 50 ),
                    OBDIVRST     => GND,
                    OBDIVHALF    => GND,
                    OBDIV0       => C ( 19 ),
                    OBDIV1       => C ( 20 ),
                    OBDIV2       => C ( 21 ),
                    OBDIV3       => C ( 22 ),
                    OBDIV4       => C ( 23 ),
                    OBMUX0       => C ( 32 ),
                    OBMUX1       => C ( 33 ),
                    OBMUX2       => C ( 34 ),
                    DLYYB0       => C ( 61 ),
                    DLYYB1       => C ( 62 ),
                    DLYYB2       => C ( 63 ),
                    DLYYB3       => C ( 64 ),
                    DLYYB4       => C ( 65 ),
                    DLYGLB0      => C ( 51 ),
                    DLYGLB1      => C ( 52 ),
                    DLYGLB2      => C ( 53 ),
                    DLYGLB3      => C ( 54 ),
                    DLYGLB4      => C ( 55 ),
                    OCDIVRST     => GND,
                    OCDIVHALF    => GND,
                    OCDIV0       => C ( 24 ),
                    OCDIV1       => C ( 25 ),
                    OCDIV2       => C ( 26 ),
                    OCDIV3       => C ( 27 ),
                    OCDIV4       => C ( 28 ),
                    OCMUX0       => C ( 35 ),
                    OCMUX1       => C ( 36 ),
                    OCMUX2       => C ( 37 ),
                    DLYYC0       => C ( 66 ),
                    DLYYC1       => C ( 67 ),
                    DLYYC2       => C ( 68 ),
                    DLYYC3       => C ( 69 ),
                    DLYYC4       => C ( 70 ),
                    DLYGLC0      => C ( 56 ),
                    DLYGLC1      => C ( 57 ),
                    DLYGLC2      => C ( 58 ),
                    DLYGLC3      => C ( 59 ),
                    DLYGLC4      => C ( 60 ),
                    FINDIV0      => C (  0 ),
                    FINDIV1      => C (  1 ),
                    FINDIV2      => C (  2 ),
                    FINDIV3      => C (  3 ),
                    FINDIV4      => C (  4 ),
                    FINDIV5      => C (  5 ),
                    FINDIV6      => C (  6 ),
                    FBDIV0       => C (  7 ),
                    FBDIV1       => C (  8 ),
                    FBDIV2       => C (  9 ),
                    FBDIV3       => C ( 10 ),
                    FBDIV4       => C ( 11 ),
                    FBDIV5       => C ( 12 ),
                    FBDIV6       => C ( 13 ),
                    FBDLY0       => C ( 40 ),
                    FBDlY1       => C ( 41 ),
                    FBDLY2       => C ( 42 ),
                    FBDLY3       => C ( 43 ),
                    FBDlY4       => C ( 44 ),
                    FBSEL0       => C ( 38 ),
                    FBSEL1       => C ( 39 ),
                    XDLYSEL      => C ( 45 ),
                    VCOSEL0      => C ( 74 ),
                    VCOSEL1      => C ( 75 ),
                    VCOSEL2      => C ( 76 ),
                    GLA          => GLA,
                    LOCK         => LOCK,
                    GLB          => GLB,
                    YB           => YB,
                    GLC          => GLC,
                    YC           => YC
                  );

  SH1: SHREG port map ( 
                    SDIN         => SDIN_ipd,
                    SCLK         => SCLK_ipd,
                    SSHIFT       => SSHIFT_ipd,
                    SUPDATE      => SUPDATE_ipd,
                    SDOUT        => SDOUT_zd,
                    SUPDATELATCH => SUPDATELATCH
                  );


  -- #########################################################
  -- # Behavior Section for timing checks
  -- #########################################################

  VITALBehavior : process ( SCLK_ipd, SSHIFT_ipd, SDIN_ipd, SUPDATE_ipd, SDOUT_zd )

     --  timing check results
     variable Tviol_SSHIFT_SCLK_posedge : X01 := '0';
     variable TmDt_SSHIFT_SCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDIN_SCLK_posedge   : X01 := '0';
     variable TmDt_SDIN_SCLK_posedge    : VitalTimingDataType := VitalTimingDataInit;

     variable Pviol_SCLK                : X01 := '0';
     variable PeriodData_SCLK           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_SUPDATE             : X01 := '0';
     variable PeriodData_SUPDATE        : VitalPeriodDataType := VitalPeriodDataInit;

     -- Output Glitch Detection Support Variables

     variable SDOUT_GlitchData          : VitalGlitchDataType;

  begin -- process VITALBehavior

  if (TimingChecksOn) then

     -- setup, hold timing check between SSHIFT and SCLK
     VitalSetupHoldCheck (
         Violation              => Tviol_SSHIFT_SCLK_posedge,
         TimingData             => TmDt_SSHIFT_SCLK_posedge,
         TestSignal             => SSHIFT_ipd,
         TestSignalName         => "SSHIFT",
         TestDelay              => 0.0 ns,
         RefSignal              => SCLK_ipd,
         RefSignalName          => "SCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_SSHIFT_SCLK_posedge_posedge,
         SetupLow               => tsetup_SSHIFT_SCLK_negedge_posedge,
         HoldHigh               => thold_SSHIFT_SCLK_posedge_posedge,
         HoldLow                => thold_SSHIFT_SCLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     -- setup, hold timing check between SDIN and SCLK
     VitalSetupHoldCheck (
         Violation              => Tviol_SDIN_SCLK_posedge,
         TimingData             => TmDt_SDIN_SCLK_posedge,
         TestSignal             => SDIN_ipd,
         TestSignalName         => "SDIN",
         TestDelay              => 0.0 ns,
         RefSignal              => SCLK_ipd,
         RefSignalName          => "SCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_SDIN_SCLK_posedge_posedge,
         SetupLow               => tsetup_SDIN_SCLK_negedge_posedge,
         HoldHigh               => thold_SDIN_SCLK_posedge_posedge,
         HoldLow                => thold_SDIN_SCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(SSHIFT_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     -- pulse width checks on SCLK 
     VitalPeriodPulseCheck (
         Violation              => Pviol_SCLK,
         PeriodData             => PeriodData_SCLK,
         TestSignal             => SCLK_ipd,
         TestSignalName         => "SCLK",
         TestDelay              => 0.0 ns,
         PulseWidthHigh         => tpw_SCLK_posedge,
         PulseWidthLow          => tpw_SCLK_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     -- pulse width checks on SUPDATE
     VitalPeriodPulseCheck (
         Violation              => Pviol_SUPDATE,
         PeriodData             => PeriodData_SUPDATE,
         TestSignal             => SUPDATE_ipd,
         TestSignalName         => "SUPDATE",
         TestDelay              => 0.0 ns,
         PulseWidthHigh         => tpw_SUPDATE_posedge,
         PulseWidthLow          => tpw_SUPDATE_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  end if;


  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

  VitalPathDelay01Z (
        OutSignal     => SDOUT,
        GlitchData    => SDOUT_GlitchData,
        OutSignalName => "SDOUT",
        OutTemp       => SDOUT_zd,
        Paths         => (0 => ( SCLK_ipd'last_event,
                                 VitalExtendToFillDelay ( tpd_SCLK_SDOUT ), TRUE )
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_DYNCCC_VITAL of DYNCCC is
   for VITAL_ACT
   end for;
end CFG_DYNCCC_VITAL;

library IEEE;
use IEEE.VITAL_Timing.all;
use IEEE.STD_LOGIC_1164.all;

-- SHREG shifts in 81 bits, but only bits 79 - 0 are included in the  
-- configuration bit string.  Bit 80 used as the RESET ENABLE.  Bits
-- 71 - 73 and 77 - 49 not used by simulation model.

-- entity declaration --
 entity DYNCCC_V2 is
   generic(
      VCOFREQUENCY      :  Real    := 0.0;
      f_CLKA_LOCK       :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

      TimingChecksOn    :  Boolean := True;
      InstancePath      :  STRING  := "*";
      Xon               :  Boolean := False;
      MsgOn             :  Boolean := True;

      tipd_CLKA         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_EXTFB        :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_POWERDOWN    :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_CLKC         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SDIN         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SCLK         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SSHIFT       :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_SUPDATE      :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
      tipd_MODE         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );

      tpd_CLKA_GLA      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLA     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLA :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLB     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLB :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_GLC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_GLC     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_GLC :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YB       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YB      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YB  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_YC       :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_EXTFB_YC      :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_POWERDOWN_YC  :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );
      tpd_CLKA_LOCK     :  VitalDelayType01 := ( 0.100 ns, 0.100 ns );

      tpd_SCLK_SDOUT    : VitalDelayType01  := ( 0.100 ns, 0.100 ns );

      tsetup_SSHIFT_SCLK_posedge_posedge : VitalDelayType := 0.000 ns;
      tsetup_SSHIFT_SCLK_negedge_posedge : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_posedge_posedge  : VitalDelayType := 0.000 ns;
      thold_SSHIFT_SCLK_negedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_SDIN_SCLK_posedge_posedge   : VitalDelayType := 0.000 ns;
      tsetup_SDIN_SCLK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_posedge_posedge    : VitalDelayType := 0.000 ns;
      thold_SDIN_SCLK_negedge_posedge    : VitalDelayType := 0.000 ns;

      tpw_SUPDATE_posedge                : VitalDelayType := 0.000 ns; 
      tpw_SUPDATE_negedge                : VitalDelayType := 0.000 ns; 
      tpw_SCLK_posedge                   : VitalDelayType := 0.000 ns;
      tpw_SCLK_negedge                   : VitalDelayType := 0.000 ns

      ); 

   port (
          CLKA         : in    std_ulogic;
          EXTFB        : in    std_ulogic;
          POWERDOWN    : in    std_ulogic;
          CLKB         : in    std_ulogic;
          CLKC         : in    std_ulogic;
          SDIN         : in    std_ulogic;
          SCLK         : in    std_ulogic;
          SSHIFT       : in    std_ulogic;
          SUPDATE      : in    std_ulogic;
          MODE         : in    std_ulogic;
          OADIV0       : in    std_ulogic;
          OADIV1       : in    std_ulogic;
          OADIV2       : in    std_ulogic;
          OADIV3       : in    std_ulogic;
          OADIV4       : in    std_ulogic;
          OAMUX0       : in    std_ulogic;
          OAMUX1       : in    std_ulogic;
          OAMUX2       : in    std_ulogic;
          DLYGLA0      : in    std_ulogic;
          DLYGLA1      : in    std_ulogic;
          DLYGLA2      : in    std_ulogic;
          DLYGLA3      : in    std_ulogic;
          DLYGLA4      : in    std_ulogic;
          OBDIV0       : in    std_ulogic;
          OBDIV1       : in    std_ulogic;
          OBDIV2       : in    std_ulogic;
          OBDIV3       : in    std_ulogic;
          OBDIV4       : in    std_ulogic;
          OBMUX0       : in    std_ulogic;
          OBMUX1       : in    std_ulogic;
          OBMUX2       : in    std_ulogic;
          DLYYB0       : in    std_ulogic;
          DLYYB1       : in    std_ulogic;
          DLYYB2       : in    std_ulogic;
          DLYYB3       : in    std_ulogic;
          DLYYB4       : in    std_ulogic;
          DLYGLB0      : in    std_ulogic;
          DLYGLB1      : in    std_ulogic;
          DLYGLB2      : in    std_ulogic;
          DLYGLB3      : in    std_ulogic;
          DLYGLB4      : in    std_ulogic;
          OCDIV0       : in    std_ulogic;
          OCDIV1       : in    std_ulogic;
          OCDIV2       : in    std_ulogic;
          OCDIV3       : in    std_ulogic;
          OCDIV4       : in    std_ulogic;
          OCMUX0       : in    std_ulogic;
          OCMUX1       : in    std_ulogic;
          OCMUX2       : in    std_ulogic;
          DLYYC0       : in    std_ulogic;
          DLYYC1       : in    std_ulogic;
          DLYYC2       : in    std_ulogic;
          DLYYC3       : in    std_ulogic;
          DLYYC4       : in    std_ulogic;
          DLYGLC0      : in    std_ulogic;
          DLYGLC1      : in    std_ulogic;
          DLYGLC2      : in    std_ulogic;
          DLYGLC3      : in    std_ulogic;
          DLYGLC4      : in    std_ulogic;
          FINDIV0      : in    std_ulogic;
          FINDIV1      : in    std_ulogic;
          FINDIV2      : in    std_ulogic;
          FINDIV3      : in    std_ulogic;
          FINDIV4      : in    std_ulogic;
          FINDIV5      : in    std_ulogic;
          FINDIV6      : in    std_ulogic;
          FBDIV0       : in    std_ulogic;
          FBDIV1       : in    std_ulogic;
          FBDIV2       : in    std_ulogic;
          FBDIV3       : in    std_ulogic;
          FBDIV4       : in    std_ulogic;
          FBDIV5       : in    std_ulogic;
          FBDIV6       : in    std_ulogic;
          FBDLY0       : in    std_ulogic;
          FBDlY1       : in    std_ulogic;
          FBDLY2       : in    std_ulogic;
          FBDLY3       : in    std_ulogic;
          FBDlY4       : in    std_ulogic;
          FBSEL0       : in    std_ulogic;
          FBSEL1       : in    std_ulogic;
          XDLYSEL      : in    std_ulogic;
          VCOSEL0      : in    std_ulogic;
          VCOSEL1      : in    std_ulogic;
          VCOSEL2      : in    std_ulogic;
          GLA          : out   std_ulogic;
          LOCK         : out   std_ulogic;
          GLB          : out   std_ulogic;
          YB           : out   std_ulogic;
          GLC          : out   std_ulogic;
          YC           : out   std_ulogic;
          SDOUT        : out   std_ulogic
        );

attribute VITAL_LEVEL0 of DYNCCC_V2 : entity is TRUE;
end DYNCCC_V2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.components.all;
use igloo.PLL_TIMING_V2;

architecture VITAL_ACT of DYNCCC_V2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal CLKA_ipd               : std_ulogic;
   signal EXTFB_ipd              : std_ulogic;
   signal POWERDOWN_ipd          : std_ulogic;
   signal CLKB_ipd               : std_ulogic;
   signal CLKC_ipd               : std_ulogic;
   signal SDIN_ipd               : std_ulogic;
   signal SCLK_ipd               : std_ulogic;
   signal SSHIFT_ipd             : std_ulogic;
   signal SUPDATE_ipd            : std_ulogic;
   signal MODE_ipd               : std_ulogic;

   signal C            : std_logic_vector ( 79 downto 0 ) := ( others => 'X' );
   signal SUPDATELATCH : std_logic_vector ( 80 downto 0 ) := ( others => 'X' );
   signal PC           : std_logic_vector ( 79 downto 0 ) := ( others => 'X' );

   -- Unused configuration bits
   signal DYNCSEL                : std_ulogic;
   signal DYNBSEL                : std_ulogic;
   signal DYNASEL                : std_ulogic;
   signal STATCSEL               : std_ulogic;
   signal STATBSEL               : std_ulogic;
   signal STATASEL               : std_ulogic;

   -- SDOUT SHREG port map
   signal SDOUT_zd               : std_ulogic;

   -- synchronisation trigger generated based on SUPDATE, MODE and SUPDATELATCH(80)
   signal DYNSYNC                : std_ulogic := '0';

   signal GND                    : std_logic  := '0';

   component PLLPRIM
     generic (
              VCOFREQUENCY          : Real;
              f_CLKA_LOCK           : Integer;
              EMULATED_SYSTEM_DELAY : Time;
              IN_DIV_DELAY          : Time;
              OUT_DIV_DELAY         : Time;
              MUX_DELAY             : Time;
              IN_DELAY_BYP1         : Time;
              BYP_MUX_DELAY         : Time;
              GL_DRVR_DELAY         : Time;
              Y_DRVR_DELAY          : Time;
              FB_MUX_DELAY          : Time;
              X_MUX_DELAY           : Time;
              FIN_LOCK_DELAY        : Time;
              LOCK_OUT_DELAY        : Time;
              PROG_INIT_DELAY       : Time;
              PROG_STEP_INCREMENT   : Time;
              BYP0_CLK_GL           : Time;
              CLKA_TO_REF_DELAY     : Time
             );
     port (
            DYNSYNC      : in    std_ulogic;
            CLKA         : in    std_ulogic;
            EXTFB        : in    std_ulogic;
            POWERDOWN    : in    std_ulogic;
            CLKB         : in    std_ulogic;
            CLKC         : in    std_ulogic;
            OADIVRST     : in    std_ulogic;
            OADIVHALF    : in    std_ulogic;
            OADIV0       : in    std_ulogic;
            OADIV1       : in    std_ulogic;
            OADIV2       : in    std_ulogic;
            OADIV3       : in    std_ulogic;
            OADIV4       : in    std_ulogic;
            OAMUX0       : in    std_ulogic;
            OAMUX1       : in    std_ulogic;
            OAMUX2       : in    std_ulogic;
            DLYGLA0      : in    std_ulogic;
            DLYGLA1      : in    std_ulogic;
            DLYGLA2      : in    std_ulogic;
            DLYGLA3      : in    std_ulogic;
            DLYGLA4      : in    std_ulogic;
            OBDIVRST     : in    std_ulogic;
            OBDIVHALF    : in    std_ulogic;
            OBDIV0       : in    std_ulogic;
            OBDIV1       : in    std_ulogic;
            OBDIV2       : in    std_ulogic;
            OBDIV3       : in    std_ulogic;
            OBDIV4       : in    std_ulogic;
            OBMUX0       : in    std_ulogic;
            OBMUX1       : in    std_ulogic;
            OBMUX2       : in    std_ulogic;
            DLYYB0       : in    std_ulogic;
            DLYYB1       : in    std_ulogic;
            DLYYB2       : in    std_ulogic;
            DLYYB3       : in    std_ulogic;
            DLYYB4       : in    std_ulogic;
            DLYGLB0      : in    std_ulogic;
            DLYGLB1      : in    std_ulogic;
            DLYGLB2      : in    std_ulogic;
            DLYGLB3      : in    std_ulogic;
            DLYGLB4      : in    std_ulogic;
            OCDIVRST     : in    std_ulogic;
            OCDIVHALF    : in    std_ulogic;
            OCDIV0       : in    std_ulogic;
            OCDIV1       : in    std_ulogic;
            OCDIV2       : in    std_ulogic;
            OCDIV3       : in    std_ulogic;
            OCDIV4       : in    std_ulogic;
            OCMUX0       : in    std_ulogic;
            OCMUX1       : in    std_ulogic;
            OCMUX2       : in    std_ulogic;
            DLYYC0       : in    std_ulogic;
            DLYYC1       : in    std_ulogic;
            DLYYC2       : in    std_ulogic;
            DLYYC3       : in    std_ulogic;
            DLYYC4       : in    std_ulogic;
            DLYGLC0      : in    std_ulogic;
            DLYGLC1      : in    std_ulogic;
            DLYGLC2      : in    std_ulogic;
            DLYGLC3      : in    std_ulogic;
            DLYGLC4      : in    std_ulogic;
            FINDIV0      : in    std_ulogic;
            FINDIV1      : in    std_ulogic;
            FINDIV2      : in    std_ulogic;
            FINDIV3      : in    std_ulogic;
            FINDIV4      : in    std_ulogic;
            FINDIV5      : in    std_ulogic;
            FINDIV6      : in    std_ulogic;
            FBDIV0       : in    std_ulogic;
            FBDIV1       : in    std_ulogic;
            FBDIV2       : in    std_ulogic;
            FBDIV3       : in    std_ulogic;
            FBDIV4       : in    std_ulogic;
            FBDIV5       : in    std_ulogic;
            FBDIV6       : in    std_ulogic;
            FBDLY0       : in    std_ulogic;
            FBDlY1       : in    std_ulogic;
            FBDLY2       : in    std_ulogic;
            FBDLY3       : in    std_ulogic;
            FBDlY4       : in    std_ulogic;
            FBSEL0       : in    std_ulogic;
            FBSEL1       : in    std_ulogic;
            XDLYSEL      : in    std_ulogic;
            VCOSEL0      : in    std_ulogic;
            VCOSEL1      : in    std_ulogic;
            VCOSEL2      : in    std_ulogic;
            GLA          : out   std_ulogic;
            LOCK         : out   std_ulogic;
            GLB          : out   std_ulogic;
            YB           : out   std_ulogic;
            GLC          : out   std_ulogic;
            YC           : out   std_ulogic
          );
     end component;

     component SHREG
       port (
              SDIN           :	in    std_ulogic;
              SCLK           :	in    std_ulogic;
              SSHIFT         :	in    std_ulogic;
              SUPDATE        :	in    std_ulogic;
              SDOUT          :	out   std_ulogic;
              SUPDATELATCH   :  out   std_logic_vector ( 80 downto 0 )
            );
     end component;
    
begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

      VitalWireDelay ( CLKA_ipd,      CLKA,      tipd_CLKA      );
      VitalWireDelay ( EXTFB_ipd,     EXTFB,     tipd_EXTFB     );
      VitalWireDelay ( POWERDOWN_ipd, POWERDOWN, tipd_POWERDOWN );
      VitalWireDelay ( CLKB_ipd,      CLKB,      tipd_CLKB      );
      VitalWireDelay ( CLKC_ipd,      CLKC,      tipd_CLKC      );
      VitalWireDelay ( SDIN_ipd,      SDIN,      tipd_SDIN      );
      VitalWireDelay ( SCLK_ipd,      SCLK,      tipd_SCLK      );
      VitalWireDelay ( SSHIFT_ipd,    SSHIFT,    tipd_SSHIFT    );
      VitalWireDelay ( SUPDATE_ipd,   SUPDATE,   tipd_SUPDATE   );
      VitalWireDelay ( MODE_ipd,      MODE,      tipd_MODE      );

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  
  PC <= 
        DYNCSEL  &
        DYNBSEL  &
        DYNASEL  &
        VCOSEL2  & 
        VCOSEL1  & 
        VCOSEL0  & 
        STATCSEL &
        STATBSEL &
        STATASEL &
        DLYYC4   &
        DLYYC3   &
        DLYYC2   &
        DLYYC1   &
        DLYYC0   &
        DLYYB4   &
        DLYYB3   &
        DLYYB2   &
        DLYYB1   &
        DLYYB0   &
        DLYGLC4  &
        DLYGLC3  &
        DLYGLC2  &
        DLYGLC1  &
        DLYGLC0  &
        DLYGLB4  &
        DLYGLB3  &
        DLYGLB2  &
        DLYGLB1  &
        DLYGLB0  &
        DLYGLA4  &
        DLYGLA3  &
        DLYGLA2  &
        DLYGLA1  &
        DLYGLA0  &
        XDLYSEL  &
        FBDLY4   &
        FBDLY3   &
        FBDLY2   &
        FBDLY1   &
        FBDLY0   &
        FBSEL1   &
        FBSEL0   &
        OCMUX2   &
        OCMUX1   &
        OCMUX0   &
        OBMUX2   &
        OBMUX1   &
        OBMUX0   &
        OAMUX2   &
        OAMUX1   &
        OAMUX0   &
        OCDIV4   &
        OCDIV3   &
        OCDIV2   &
        OCDIV1   &
        OCDIV0   &
        OBDIV4   &
        OBDIV3   &
        OBDIV2   &
        OBDIV1   &
        OBDIV0   &
        OADIV4   &
        OADIV3   &
        OADIV2   &
        OADIV1   &
        OADIV0   &
        FBDIV6   &
        FBDIV5   &
        FBDIV4   &
        FBDIV3   &
        FBDIV2   &
        FBDIV1   &
        FBDIV0   &
        FINDIV6  &
        FINDIV5  &
        FINDIV4  &
        FINDIV3  &
        FINDIV2  &
        FINDIV1  &
        FINDIV0  ;

  C <= SUPDATELATCH ( 79 downto 0 ) when ( TO_X01 ( MODE_ipd ) = '1' ) else
       PC ( 79 downto 0 ) when ( TO_X01 ( MODE_ipd ) = '0' ) else
       "XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX";

  -- logic for generating DYNSYNC

  latch_mode_reset : process ( SUPDATE_ipd )

    variable RESETENA_latched : std_ulogic;

  begin

    if ( TO_X01 ( SUPDATE_ipd ) = '1' ) then
      if ( TO_X01( MODE_ipd ) = '1' and TO_X01( RESETENA_latched ) = '1' ) then
        DYNSYNC <= '1'; 
      end if;
    elsif ( TO_X01 ( SUPDATE_ipd ) = '0' ) then
      DYNSYNC <= '0';
      RESETENA_latched := SUPDATELATCH ( 80 );
    end if;

  end process;


  P1: PLLPRIM 
      generic map (
                    VCOFREQUENCY          => VCOFREQUENCY,
                    f_CLKA_LOCK           => f_CLKA_LOCK,
                    EMULATED_SYSTEM_DELAY => PLL_TIMING_V2.EMULATED_SYSTEM_DELAY,
                    IN_DIV_DELAY          => PLL_TIMING_V2.IN_DIV_DELAY,
                    OUT_DIV_DELAY         => PLL_TIMING_V2.OUT_DIV_DELAY,
                    MUX_DELAY             => PLL_TIMING_V2.MUX_DELAY,
                    IN_DELAY_BYP1         => PLL_TIMING_V2.IN_DELAY_BYP1,
                    BYP_MUX_DELAY         => PLL_TIMING_V2.BYP_MUX_DELAY,
                    GL_DRVR_DELAY         => PLL_TIMING_V2.GL_DRVR_DELAY,
                    Y_DRVR_DELAY          => PLL_TIMING_V2.Y_DRVR_DELAY,
                    FB_MUX_DELAY          => PLL_TIMING_V2.FB_MUX_DELAY,
                    X_MUX_DELAY           => PLL_TIMING_V2.X_MUX_DELAY,
                    FIN_LOCK_DELAY        => PLL_TIMING_V2.FIN_LOCK_DELAY,
                    LOCK_OUT_DELAY        => PLL_TIMING_V2.LOCK_OUT_DELAY,
                    PROG_INIT_DELAY       => PLL_TIMING_V2.PROG_INIT_DELAY,
                    PROG_STEP_INCREMENT   => PLL_TIMING_V2.PROG_STEP_INCREMENT,
                    BYP0_CLK_GL           => PLL_TIMING_V2.BYP0_CLK_GL,
                    CLKA_TO_REF_DELAY     => PLL_TIMING_V2.CLKA_TO_REF_DELAY
                  )
      port map    ( 
                    DYNSYNC      => DYNSYNC,
                    CLKA         => CLKA_ipd,
                    EXTFB        => EXTFB_ipd,
                    POWERDOWN    => POWERDOWN_ipd,
                    CLKB         => CLKB_ipd,
                    CLKC         => CLKC_ipd,
                    OADIVRST     => GND,
                    OADIVHALF    => GND,
                    OADIV0       => C ( 14 ),
                    OADIV1       => C ( 15 ),
                    OADIV2       => C ( 16 ),
                    OADIV3       => C ( 17 ),
                    OADIV4       => C ( 18 ),
                    OAMUX0       => C ( 29 ),
                    OAMUX1       => C ( 30 ),
                    OAMUX2       => C ( 31 ),
                    DLYGLA0      => C ( 46 ),
                    DLYGLA1      => C ( 47 ),
                    DLYGLA2      => C ( 48 ),
                    DLYGLA3      => C ( 49 ),
                    DLYGLA4      => C ( 50 ),
                    OBDIVRST     => GND,
                    OBDIVHALF    => GND,
                    OBDIV0       => C ( 19 ),
                    OBDIV1       => C ( 20 ),
                    OBDIV2       => C ( 21 ),
                    OBDIV3       => C ( 22 ),
                    OBDIV4       => C ( 23 ),
                    OBMUX0       => C ( 32 ),
                    OBMUX1       => C ( 33 ),
                    OBMUX2       => C ( 34 ),
                    DLYYB0       => C ( 61 ),
                    DLYYB1       => C ( 62 ),
                    DLYYB2       => C ( 63 ),
                    DLYYB3       => C ( 64 ),
                    DLYYB4       => C ( 65 ),
                    DLYGLB0      => C ( 51 ),
                    DLYGLB1      => C ( 52 ),
                    DLYGLB2      => C ( 53 ),
                    DLYGLB3      => C ( 54 ),
                    DLYGLB4      => C ( 55 ),
                    OCDIVRST     => GND,
                    OCDIVHALF    => GND,
                    OCDIV0       => C ( 24 ),
                    OCDIV1       => C ( 25 ),
                    OCDIV2       => C ( 26 ),
                    OCDIV3       => C ( 27 ),
                    OCDIV4       => C ( 28 ),
                    OCMUX0       => C ( 35 ),
                    OCMUX1       => C ( 36 ),
                    OCMUX2       => C ( 37 ),
                    DLYYC0       => C ( 66 ),
                    DLYYC1       => C ( 67 ),
                    DLYYC2       => C ( 68 ),
                    DLYYC3       => C ( 69 ),
                    DLYYC4       => C ( 70 ),
                    DLYGLC0      => C ( 56 ),
                    DLYGLC1      => C ( 57 ),
                    DLYGLC2      => C ( 58 ),
                    DLYGLC3      => C ( 59 ),
                    DLYGLC4      => C ( 60 ),
                    FINDIV0      => C (  0 ),
                    FINDIV1      => C (  1 ),
                    FINDIV2      => C (  2 ),
                    FINDIV3      => C (  3 ),
                    FINDIV4      => C (  4 ),
                    FINDIV5      => C (  5 ),
                    FINDIV6      => C (  6 ),
                    FBDIV0       => C (  7 ),
                    FBDIV1       => C (  8 ),
                    FBDIV2       => C (  9 ),
                    FBDIV3       => C ( 10 ),
                    FBDIV4       => C ( 11 ),
                    FBDIV5       => C ( 12 ),
                    FBDIV6       => C ( 13 ),
                    FBDLY0       => C ( 40 ),
                    FBDlY1       => C ( 41 ),
                    FBDLY2       => C ( 42 ),
                    FBDLY3       => C ( 43 ),
                    FBDlY4       => C ( 44 ),
                    FBSEL0       => C ( 38 ),
                    FBSEL1       => C ( 39 ),
                    XDLYSEL      => C ( 45 ),
                    VCOSEL0      => C ( 74 ),
                    VCOSEL1      => C ( 75 ),
                    VCOSEL2      => C ( 76 ),
                    GLA          => GLA,
                    LOCK         => LOCK,
                    GLB          => GLB,
                    YB           => YB,
                    GLC          => GLC,
                    YC           => YC
                  );

  SH1: SHREG port map ( 
                    SDIN         => SDIN_ipd,
                    SCLK         => SCLK_ipd,
                    SSHIFT       => SSHIFT_ipd,
                    SUPDATE      => SUPDATE_ipd,
                    SDOUT        => SDOUT_zd,
                    SUPDATELATCH => SUPDATELATCH
                  );


  -- #########################################################
  -- # Behavior Section for timing checks
  -- #########################################################

  VITALBehavior : process ( SCLK_ipd, SSHIFT_ipd, SDIN_ipd, SUPDATE_ipd, SDOUT_zd )

     --  timing check results
     variable Tviol_SSHIFT_SCLK_posedge : X01 := '0';
     variable TmDt_SSHIFT_SCLK_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_SDIN_SCLK_posedge   : X01 := '0';
     variable TmDt_SDIN_SCLK_posedge    : VitalTimingDataType := VitalTimingDataInit;

     variable Pviol_SCLK                : X01 := '0';
     variable PeriodData_SCLK           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_SUPDATE             : X01 := '0';
     variable PeriodData_SUPDATE        : VitalPeriodDataType := VitalPeriodDataInit;

     -- Output Glitch Detection Support Variables

     variable SDOUT_GlitchData          : VitalGlitchDataType;

  begin -- process VITALBehavior

  if (TimingChecksOn) then

     -- setup, hold timing check between SSHIFT and SCLK
     VitalSetupHoldCheck (
         Violation              => Tviol_SSHIFT_SCLK_posedge,
         TimingData             => TmDt_SSHIFT_SCLK_posedge,
         TestSignal             => SSHIFT_ipd,
         TestSignalName         => "SSHIFT",
         TestDelay              => 0.0 ns,
         RefSignal              => SCLK_ipd,
         RefSignalName          => "SCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_SSHIFT_SCLK_posedge_posedge,
         SetupLow               => tsetup_SSHIFT_SCLK_negedge_posedge,
         HoldHigh               => thold_SSHIFT_SCLK_posedge_posedge,
         HoldLow                => thold_SSHIFT_SCLK_negedge_posedge,
         CheckEnabled           => TRUE,
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     -- setup, hold timing check between SDIN and SCLK
     VitalSetupHoldCheck (
         Violation              => Tviol_SDIN_SCLK_posedge,
         TimingData             => TmDt_SDIN_SCLK_posedge,
         TestSignal             => SDIN_ipd,
         TestSignalName         => "SDIN",
         TestDelay              => 0.0 ns,
         RefSignal              => SCLK_ipd,
         RefSignalName          => "SCLK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_SDIN_SCLK_posedge_posedge,
         SetupLow               => tsetup_SDIN_SCLK_negedge_posedge,
         HoldHigh               => thold_SDIN_SCLK_posedge_posedge,
         HoldLow                => thold_SDIN_SCLK_negedge_posedge,
         CheckEnabled           => (TO_X01(SSHIFT_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     -- pulse width checks on SCLK 
     VitalPeriodPulseCheck (
         Violation              => Pviol_SCLK,
         PeriodData             => PeriodData_SCLK,
         TestSignal             => SCLK_ipd,
         TestSignalName         => "SCLK",
         TestDelay              => 0.0 ns,
         PulseWidthHigh         => tpw_SCLK_posedge,
         PulseWidthLow          => tpw_SCLK_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

     -- pulse width checks on SUPDATE
     VitalPeriodPulseCheck (
         Violation              => Pviol_SUPDATE,
         PeriodData             => PeriodData_SUPDATE,
         TestSignal             => SUPDATE_ipd,
         TestSignalName         => "SUPDATE",
         TestDelay              => 0.0 ns,
         PulseWidthHigh         => tpw_SUPDATE_posedge,
         PulseWidthLow          => tpw_SUPDATE_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/DYNCCC",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  end if;


  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

  VitalPathDelay01Z (
        OutSignal     => SDOUT,
        GlitchData    => SDOUT_GlitchData,
        OutSignalName => "SDOUT",
        OutTemp       => SDOUT_zd,
        Paths         => (0 => ( SCLK_ipd'last_event,
                                 VitalExtendToFillDelay ( tpd_SCLK_SDOUT ), TRUE )
                         ),
        DefaultDelay  => VitalZeroDelay01Z,
        Mode          => Onevent,
        XON           => Xon,
        MsgOn         => MsgOn,
        MsgSeverity   => WARNING
        );

  end process VITALBehavior;

end VITAL_ACT;

configuration CFG_DYNCCC_V2_VITAL of DYNCCC_V2 is
   for VITAL_ACT
   end for;
end CFG_DYNCCC_V2_VITAL;

----- CELL UJTAG -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity UJTAG is
   generic(
      TimingChecksOn : Boolean := True;
      InstancePath   : STRING  := "*";
      Xon            : Boolean := False;
      MsgOn          : Boolean := True;

      tipd_UTDO        : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TMS         : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TDI         : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TCK         : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TRSTB       : VitalDelayType01 := (0.0 ns, 0.0 ns);

      tpd_TCK_UIREG0   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG1   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG2   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG3   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG4   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG5   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG6   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UIREG7   : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TCK_URSTB    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRSH    : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRCAP   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRUPD   : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TCK_UDRCK    : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TCK_TDO      : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TRSTB_UIREG0 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG1 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG2 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG3 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG4 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG5 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG6 : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UIREG7 : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TRSTB_URSTB  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UDRSH  : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UDRCAP : VitalDelayType01 := (0.100 ns, 0.100 ns);
      tpd_TRSTB_UDRUPD : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TRSTB_TDO    : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tpd_TDI_UTDI     : VitalDelayType01 := (0.100 ns, 0.100 ns);

      tsetup_TDI_TCK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_TDI_TCK_negedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_TMS_TCK_posedge_posedge  : VitalDelayType := 0.000 ns;
      tsetup_TMS_TCK_negedge_posedge  : VitalDelayType := 0.000 ns;

      tsetup_UTDO_TCK_posedge_negedge : VitalDelayType := 0.000 ns;
      tsetup_UTDO_TCK_negedge_negedge : VitalDelayType := 0.000 ns;

      thold_TDI_TCK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_TDI_TCK_negedge_posedge   : VitalDelayType := 0.000 ns;
      thold_TMS_TCK_posedge_posedge   : VitalDelayType := 0.000 ns;
      thold_TMS_TCK_negedge_posedge   : VitalDelayType := 0.000 ns;

      thold_UTDO_TCK_posedge_negedge  : VitalDelayType := 0.000 ns;
      thold_UTDO_TCK_negedge_negedge  : VitalDelayType := 0.000 ns;

      trecovery_TRSTB_TCK_posedge_posedge : VitalDelayType := 0.000 ns;
      thold_TRSTB_TCK_posedge_posedge     : VitalDelayType := 0.000 ns;

      tpw_TCK_posedge   : VitalDelayType := 0.000 ns;
      tpw_TCK_negedge   : VitalDelayType := 0.000 ns;
      tpw_TRSTB_negedge : VitalDelayType := 0.000 ns

     );

   port(
      UTDO           :	in    STD_ULOGIC; 
      TMS            :	in    STD_ULOGIC;
      TDI            :	in    STD_ULOGIC;  
      TCK            :	in    STD_ULOGIC;
      TRSTB          :	in    STD_ULOGIC; 
      UIREG0         :  out   STD_ULOGIC;
      UIREG1         :  out   STD_ULOGIC;
      UIREG2         :  out   STD_ULOGIC;
      UIREG3         :  out   STD_ULOGIC;
      UIREG4         :  out   STD_ULOGIC;
      UIREG5         :  out   STD_ULOGIC;
      UIREG6         :  out   STD_ULOGIC;
      UIREG7         :  out   STD_ULOGIC;
      UTDI           :  out   STD_ULOGIC;
      URSTB          :  out   STD_ULOGIC;
      UDRCK          :  out   STD_ULOGIC;
      UDRCAP         :  out   STD_ULOGIC;
      UDRSH          :  out   STD_ULOGIC;
      UDRUPD         :  out   STD_ULOGIC;
      TDO            :  out   STD_ULOGIC);            

  attribute VITAL_LEVEL0 of UJTAG : entity is TRUE;
end UJTAG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of UJTAG is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL UTDO_ipd          : STD_ULOGIC := 'X';
   SIGNAL TMS_ipd           : STD_ULOGIC := 'X';
   SIGNAL TDI_ipd           : STD_ULOGIC := 'X';
   SIGNAL TCK_ipd           : STD_ULOGIC := 'X';
   SIGNAL TRSTB_ipd         : STD_ULOGIC := 'X';

   SIGNAL SHREG             : std_logic_vector(7 downto 0) := "XXXXXXXX";
   SIGNAL IR                : std_logic_vector(7 downto 0);

   type state_type is (Test_Logic_Reset,
                       Run_Test_Idle,
                       Select_DR,
                       Capture_DR,
                       Shift_DR,
                       Exit1_DR,
                       Pause_DR,
                       Exit2_DR,
                       Update_DR,
                       Select_IR,
                       Capture_IR,
                       Shift_IR,
                       Exit1_IR,
                       Pause_IR,
                       Exit2_IR,
                       Update_IR,
                       Unknown
                      );

   SIGNAL STATE : state_type := Unknown;

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

     VitalWireDelay (UTDO_ipd, UTDO, tipd_UTDO);
     VitalWireDelay (TMS_ipd, TMS, tipd_TMS);
     VitalWireDelay (TDI_ipd, TDI, tipd_TDI);
     VitalWireDelay (TCK_ipd, TCK, tipd_TCK);
     VitalWireDelay (TRSTB_ipd, TRSTB, tipd_TRSTB);

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  OUTPUTS1 : process (TCK_ipd, TRSTB_ipd, TMS_ipd, TDI_ipd, UTDO_ipd )

  --  Timing Check Results
  variable Tviol_TDI_TCK_posedge  : X01 := '0';
  variable TmDt_TDI_TCK_posedge   : VitalTimingDataType := VitalTimingDataInit;
  variable Tviol_TMS_TCK_posedge  : X01 := '0';
  variable TmDt_TMS_TCK_posedge   : VitalTimingDataType := VitalTimingDataInit;
  variable Tviol_UTDO_TCK_negedge : X01 := '0';
  variable TmDt_UTDO_TCK_negedge  : VitalTimingDataType := VitalTimingDataInit;

  variable Pviol_TCK                : X01 := '0';
  variable PeriodData_TCK           : VitalPeriodDataType := VitalPeriodDataInit;
  variable Tviol_TRSTB_TCK_posedge  : X01 := '0';
  variable Tmkr_TRSTB_TCK_posedge   : VitalTimingDataType := VitalTimingDataInit;
  variable Pviol_TRSTB              : X01 := '0';
  variable PeriodData_TRSTB         : VitalPeriodDataType := VitalPeriodDataInit;

  -- functional Results
  variable UDRUPD_zd : std_ulogic;
  variable UDRSH_zd  : std_ulogic;
  variable UDRCAP_zd : std_ulogic;
  variable URSTB_zd  : std_ulogic;

  -- Output Glitch Detection Support Variables
  variable UDRUPD_GlitchData : VitalGlitchDataType;
  variable UDRSH_GlitchData  : VitalGlitchDataType;
  variable UDRCAP_GlitchData : VitalGlitchDataType;
  variable URSTB_GlitchData  : VitalGlitchDataType;

  begin

  if (TimingChecksOn) then
  ---------------------------------------------------------
  -- # Timing Check Section                              --
  ---------------------------------------------------------

  -- recovery/ removal check for TCK to TRSTB signal
    VitalRecoveryRemovalCheck   (
         Violation              => Tviol_TRSTB_TCK_posedge,
         TimingData             => Tmkr_TRSTB_TCK_posedge,
         TestSignal             => TRSTB_ipd,
         TestSignalName         => "TRSTB",
         TestDelay              => 0 ns,
         RefSignal              => TCK_ipd,
         RefSignalName          => "TCK",
         RefDelay               => 0 ns,
         Recovery               => trecovery_TRSTB_TCK_posedge_posedge,
         Removal                => thold_TRSTB_TCK_posedge_posedge,
         ActiveLow              => TRUE,
         CheckEnabled           => TRUE,
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/UJTAG",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING);

  -- setup / hold TDI to TCK
    VitalSetupHoldCheck (
         Violation              => Tviol_TDI_TCK_posedge,
         TimingData             => TmDt_TDI_TCK_posedge,
         TestSignal             => TDI_ipd,
         TestSignalName         => "TDI",
         TestDelay              => 0.0 ns,
         RefSignal              => TCK_ipd,
         RefSignalName          => "TCK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_TDI_TCK_posedge_posedge,
         SetupLow               => tsetup_TDI_TCK_negedge_posedge,
         HoldHigh               => thold_TDI_TCK_posedge_posedge,
         HoldLow                => thold_TDI_TCK_negedge_posedge,
         CheckEnabled           => (TO_X01(TRSTB_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/UJTAG",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- setup / hold TMS to TCK
    VitalSetupHoldCheck (
         Violation              => Tviol_TMS_TCK_posedge,
         TimingData             => TmDt_TMS_TCK_posedge,
         TestSignal             => TMS_ipd,
         TestSignalName         => "TMS",
         TestDelay              => 0.0 ns,
         RefSignal              => TCK_ipd,
         RefSignalName          => "TCK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_TMS_TCK_posedge_posedge,
         SetupLow               => tsetup_TMS_TCK_negedge_posedge,
         HoldHigh               => thold_TMS_TCK_posedge_posedge,
         HoldLow                => thold_TMS_TCK_negedge_posedge,
         CheckEnabled           => (TO_X01(TRSTB_ipd) = '1'),
         RefTransition          => '/',
         HeaderMsg              => InstancePath & "/UJTAG",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  -- setup / hold UTDO to TCK
    VitalSetupHoldCheck (
         Violation              => Tviol_UTDO_TCK_negedge,
         TimingData             => TmDt_UTDO_TCK_negedge,
         TestSignal             => UTDO_ipd,
         TestSignalName         => "UTDO",
         TestDelay              => 0.0 ns,
         RefSignal              => TCK_ipd,
         RefSignalName          => "TCK",
         RefDelay               => 0.0 ns,
         SetupHigh              => tsetup_UTDO_TCK_posedge_negedge,
         SetupLow               => tsetup_UTDO_TCK_negedge_negedge,
         HoldHigh               => thold_UTDO_TCK_posedge_negedge,
         HoldLow                => thold_UTDO_TCK_negedge_negedge,
         CheckEnabled           => (TO_X01(TRSTB_ipd) = '1'),
         RefTransition          => '\',
         HeaderMsg              => InstancePath & "/UJTAG",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  --  Period of TCK
    VitalPeriodPulseCheck (
         Violation              => Pviol_TCK,
         PeriodData             => PeriodData_TCK,
         TestSignal             => TCK_ipd,
         TestSignalName         => "TCK",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => tpw_TCK_posedge,
         PulseWidthLow          => tpw_TCK_negedge,
         CheckEnabled           => (TO_X01(TRSTB_ipd) = '1'),
         HeaderMsg              => InstancePath & "/UJTAG",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

  --  Period of TRSTB
    VitalPeriodPulseCheck (
         Violation              => Pviol_TRSTB,
         PeriodData             => PeriodData_TRSTB,
         TestSignal             => TRSTB_ipd,
         TestSignalName         => "TRSTB",
         TestDelay              => 0.0 ns,
         Period                 => 0.0 ns,
         PulseWidthHigh         => 0.0 ns,
         PulseWidthLow          => tpw_TRSTB_negedge,
         CheckEnabled           => TRUE,
         HeaderMsg              => InstancePath & "/UJTAG",
         Xon                    => Xon,
         MsgOn                  => MsgOn,
         MsgSeverity            => WARNING
         );

   end if;

    if ((TRSTB_ipd'event) and (TO_X01(TRSTB_ipd) = '0')) then
                UDRUPD_zd := '0';
                UDRSH_zd  := '0';
                UDRCAP_zd := '0';
                URSTB_zd  := '0';
  
    elsif ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '0')) then
      if (STATE = Unknown) then
        UDRUPD_zd := 'X';
        UDRSH_zd  := 'X';
        UDRCAP_zd := 'X';
        URSTB_zd  := 'X';
      else
        if (STATE = Update_DR) then
          UDRUPD_zd := '1';
        else
          UDRUPD_zd := '0';
        end if;
    
        if (STATE = Shift_DR) then
          UDRSH_zd  := '1';
        else
          UDRSH_zd  := '0';
        end if;

        if (STATE = Capture_DR) then
          UDRCAP_zd := '1';
        else
          UDRCAP_zd := '0';
        end if;
        
        if(STATE /= Test_Logic_Reset) then
          URSTB_zd  := '1';
        else
          URSTB_zd  := '0';
        end if;
      end if;
    end if;

  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

  VitalPathDelay01Z (
    OutSignal     => UDRUPD,
    GlitchData    => UDRUPD_GlitchData,
    OutSignalName => "UDRUPD",
    OutTemp       => UDRUPD_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UDRUPD), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UDRUPD), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UDRSH,
    GlitchData    => UDRSH_GlitchData,
    OutSignalName => "UDRSH",
    OutTemp       => UDRSH_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UDRSH), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UDRSH), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UDRCAP,
    GlitchData    => UDRCAP_GlitchData,
    OutSignalName => "UDRCAP",
    OutTemp       => UDRCAP_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UDRCAP), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UDRCAP), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => URSTB,
    GlitchData    => URSTB_GlitchData,
    OutSignalName => "URSTB",
    OutTemp       => URSTB_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_URSTB), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_URSTB), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  end process OUTPUTS1;

  STATES: process (TCK_ipd, TRSTB_ipd)
  begin
    if ((TRSTB_ipd'event) and (TO_X01(TRSTB_ipd) = '0')) then
       STATE <= Test_Logic_Reset;
    elsif ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '1')) then
       case STATE is
         when Test_Logic_Reset       => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Test_Logic_Reset;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Run_Test_Idle;
                                        end if;
         when Run_Test_Idle          => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Select_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Run_Test_Idle;
                                        end if;
         when Select_DR              => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Select_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Capture_DR;
                                        end if;
         when Capture_DR | Shift_DR  => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Exit1_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_DR;
                                        end if;
         when Exit1_DR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_DR;
                                        end if;
         when Pause_DR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Exit2_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_DR;
                                        end if;
         when Exit2_DR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_DR;
                                        end if;
         when  Select_IR             => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Test_Logic_Reset;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Capture_IR;
                                        end if;
         when Capture_IR | Shift_IR  => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Exit1_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_IR;
                                        end if;
         when Exit1_IR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_IR;
                                        end if;
         when Pause_IR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <=  Exit2_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_IR;
                                        end if;
         when Exit2_IR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_IR;
                                        end if;
         when Update_DR | Update_IR  => if (TO_X01(TMS_ipd)= '1') then
                                          STATE <= Select_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Run_Test_Idle;
                                        end if;
         when Unknown                => STATE <= Unknown;
       end case;
    end if;
  end process STATES;

  CLOCK_SHREG: process(TCK_ipd)
  begin
    if ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '1')) then
      case STATE is
        when Capture_IR  => SHREG <=  "XXXXXX01";
        when Capture_DR  => SHREG <=  "00000000";
        when Shift_IR | Shift_DR  => SHREG <= TDI_ipd & SHREG(7) & SHREG(6) & SHREG(5) 
                                              & SHREG(4) & SHREG(3) & SHREG(2) & SHREG(1);
    
        when others   => SHREG <= SHREG;  
      end case;
    end if;
  end process CLOCK_SHREG;


  OUTPUTS2: process(TCK_ipd, TRSTB_ipd)

  -- functional Results

  variable TDO_zd    : std_ulogic;
  variable UIREG0_zd : std_ulogic;
  variable UIREG1_zd : std_ulogic;
  variable UIREG2_zd : std_ulogic;
  variable UIREG3_zd : std_ulogic;
  variable UIREG4_zd : std_ulogic;
  variable UIREG5_zd : std_ulogic;
  variable UIREG6_zd : std_ulogic;
  variable UIREG7_zd : std_ulogic;
  variable UDRCK_zd  : std_ulogic;

  -- Output Glitch Detection Support Variables
  variable TDO_GlitchData    : VitalGlitchDataType;
  variable UIREG0_GlitchData : VitalGlitchDataType;
  variable UIREG1_GlitchData : VitalGlitchDataType;
  variable UIREG2_GlitchData : VitalGlitchDataType;
  variable UIREG3_GlitchData : VitalGlitchDataType;
  variable UIREG4_GlitchData : VitalGlitchDataType;
  variable UIREG5_GlitchData : VitalGlitchDataType;
  variable UIREG6_GlitchData : VitalGlitchDataType;
  variable UIREG7_GlitchData : VitalGlitchDataType;
  variable UDRCK_GlitchData  : VitalGlitchDataType;

  begin
    UDRCK_zd := TCK_ipd;
    if ((TRSTB_ipd'event) and (TO_X01(TRSTB_ipd) = '0')) then
      IR        <= "11111111"; -- Bypass
      UIREG0_zd := '1'; 
      UIREG1_zd := '1';
      UIREG2_zd := '1';
      UIREG3_zd := '1';
      UIREG4_zd := '1';
      UIREG5_zd := '1';
      UIREG6_zd := '1';
      UIREG7_zd := '1';
      TDO_zd    := 'Z';
    elsif ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '0')) then
      if (STATE = Shift_IR) then
        TDO_zd := SHREG(0);
      elsif (STATE = Shift_DR) then
        if (IR(7) = '0' and (IR(6) = '1' or IR(5) = '1' or IR(4) = '1')) then
          TDO_zd := UTDO;
        else
          TDO_zd := SHREG(7);
        end if;
      elsif (STATE = Update_IR) then
        TDO_zd    := 'Z';
        IR        <= SHREG;
        UIREG0_zd := SHREG(0);
        UIREG1_zd := SHREG(1);
        UIREG2_zd := SHREG(2);
        UIREG3_zd := SHREG(3);
        UIREG4_zd := SHREG(4);
        UIREG5_zd := SHREG(5);
        UIREG6_zd := SHREG(6);
        UIREG7_zd := SHREG(7);
      else
        TDO_zd := 'Z';
      end if;
    end if;

  -- #########################################################
  -- # Path Delay Section
  -- #########################################################

  VitalPathDelay01Z (
    OutSignal     => TDO,
    GlitchData    => TDO_GlitchData,
    OutSignalName => "TDO",
    OutTemp       => TDO_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_TDO), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_TDO), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG0,
    GlitchData    => UIREG0_GlitchData,
    OutSignalName => "UIREG0",
    OutTemp       => UIREG0_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG0), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG0), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG1,
    GlitchData    => UIREG1_GlitchData,
    OutSignalName => "UIREG1",
    OutTemp       => UIREG1_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG1), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG1), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG2,
    GlitchData    => UIREG2_GlitchData,
    OutSignalName => "UIREG2",
    OutTemp       => UIREG2_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG2), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG2), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG3,
    GlitchData    => UIREG3_GlitchData,
    OutSignalName => "UIREG3",
    OutTemp       => UIREG3_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG3), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG3), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG4,
    GlitchData    => UIREG4_GlitchData,
    OutSignalName => "UIREG4",
    OutTemp       => UIREG4_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG4), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG4), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG5,
    GlitchData    => UIREG5_GlitchData,
    OutSignalName => "UIREG5",
    OutTemp       => UIREG5_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG5), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG5), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG6,
    GlitchData    => UIREG6_GlitchData,
    OutSignalName => "UIREG6",
    OutTemp       => UIREG6_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG6), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG6), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UIREG7,
    GlitchData    => UIREG7_GlitchData,
    OutSignalName => "UIREG7",
    OutTemp       => UIREG7_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UIREG7), TRUE),
                      1 => (TRSTB_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TRSTB_UIREG7), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );

  VitalPathDelay01Z (
    OutSignal     => UDRCK,
    GlitchData    => UDRCK_GlitchData,
    OutSignalName => "UDRCK",
    OutTemp       => UDRCK_zd,
    Paths         => (0 => (TCK_ipd'last_event,
                            VitalExtendToFillDelay(tpd_TCK_UDRCK), TRUE)
                     ),
    DefaultDelay  => VitalZeroDelay01Z,
    Mode          => Onevent,
    XON           => Xon,
    MsgOn         => MsgOn,
    MsgSeverity   => WARNING
  );
  
  end process OUTPUTS2;

--  OUTPUTS3: process(IR)
--  begin
--    UIREG7 <= IR(7);
--    UIREG6 <= IR(6);
--    UIREG5 <= IR(5);
--    UIREG4 <= IR(4);
--    UIREG3 <= IR(3);
--    UIREG2 <= IR(2);
--    UIREG1 <= IR(1);
--    UIREG0 <= IR(0);
--  end process OUTPUTS3;

  OUTPUTS4: process(TDI_ipd)

  -- functional Results
  variable UTDI_zd    : std_ulogic;
                            
  -- Output Glitch Detection Support Variables
  variable UTDI_GlitchData    : VitalGlitchDataType;

  begin

    UTDI_zd := TDI_ipd;

    VitalPathDelay01Z (
      OutSignal     => UTDI,
      GlitchData    => UTDI_GlitchData,
      OutSignalName => "UTDI",
      OutTemp       => UTDI_zd,
      Paths         => (0 => (TDI_ipd'last_event,
                              VitalExtendToFillDelay(tpd_TDI_UTDI), TRUE)
                       ),
      DefaultDelay  => VitalZeroDelay01Z,
      Mode          => Onevent,
      XON           => Xon,
      MsgOn         => MsgOn,
      MsgSeverity   => WARNING
    );

  end process;

-- UTDI <= TDI_ipd;

--  OUTPUTS5: process(TCK_ipd)
--  begin
--    UDRCK <= TCK_ipd;
--  end process;

-- UDRCK_zd <= TCK_ipd;

--  OUTPUTS6: process(STATE)
--  begin
--    if (STATE = Unknown) then
--      URSTB <= 'X';
--    elsif (STATE = Test_Logic_Reset) then
--      URSTB <= '0';
--    else
--      URSTB <= '1';
--   end if;
--  end process;


end VITAL_ACT;

configuration CFG_UJTAG_VITAL of UJTAG is
  for VITAL_ACT
  end for;
end CFG_UJTAG_VITAL;


 ---- CELL SIMBUF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;

 ---- entity declaration ----
 entity SIMBUF is

    port(
		D		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end SIMBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library igloo;
use igloo.VTABLES.all;

architecture VITAL_ACT of SIMBUF is
begin
        PAD <= TO_X01(D);
end VITAL_ACT;

 configuration CFG_SIMBUF_VITAL of SIMBUF is 
    for VITAL_ACT
    end for;
 end CFG_SIMBUF_VITAL;
--***************************************************************************

--***************************************************************************
-- Detailed Revision History:
--
-- Version  Date(MM/DD/YY)   Submitter              Description
--
-- 1.0      10/8/09         Kiran Yerribandi     First Version.
--------------------------------------------------------------------
-- CELL NAME : PLL_SDF
---------------------------------------------------------------------

--  PLL_SDF and PLL_DLY_SDF macros are used to model backannotated pll model.
--  In the backannotated netlist PLL is split up into two macros PLL_SDF and
--  PLL_DLY_SDF. PLL_SDF macro has all the functionality and PLL_DLY_SDF
--  modules all the delays.
-- PLL_SDF macro doesn;t have any delays in it.
--     #########################################################
--     #                    PLLBA                              #   
--     #                                                       #
--     #     ----------               -----------              #
--     #    |          |             |           |             #
--     #    |          |-----------> |           |             #
--     #    |PLL_SDF   |             |PLL_DLY_SDF|             #
--     #    |          |             |           |             #
--     #    |          |             |           |             #
--     #    |          |             |           |---          #
--     #  --|          |             |           |   |         #
--     #  |  ----------               -----------    |         #
--     #  |                                          |         #
--     #   -------------------------------------------         #
--     #                                                       #
--     #########################################################

library IEEE;
use IEEE.std_logic_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity PLL_SDF is
  generic (
    VCOFREQUENCY       :  Real    := 0.0;
    f_CLKA_LOCK        :  Integer := 3; -- Number of CLKA pulses after which LOCK is raised

    TimingChecksOn     :  Boolean          := True;
    InstancePath       :  String           := "*";
    Xon                :  Boolean          := False;
    MsgOn              :  Boolean          := True;
    tipd_CLKA          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_EXTFB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_INTFB         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tipd_POWERDOWN     :  VitalDelayType01 := ( 0.000 ns, 0.000 ns )
   );

  port (
    CLKA         : in    std_ulogic;
    EXTFB        : in    std_ulogic;
    INTFB        : in    std_ulogic;
    POWERDOWN    : in    std_ulogic;
    OADIV0       : in    std_ulogic;
    OADIV1       : in    std_ulogic;
    OADIV2       : in    std_ulogic;
    OADIV3       : in    std_ulogic;
    OADIV4       : in    std_ulogic;
    OAMUX0       : in    std_ulogic;
    OAMUX1       : in    std_ulogic;
    OAMUX2       : in    std_ulogic;
    DLYGLA0      : in    std_ulogic;
    DLYGLA1      : in    std_ulogic;
    DLYGLA2      : in    std_ulogic;
    DLYGLA3      : in    std_ulogic;
    DLYGLA4      : in    std_ulogic;
    OBDIV0       : in    std_ulogic;
    OBDIV1       : in    std_ulogic;
    OBDIV2       : in    std_ulogic;
    OBDIV3       : in    std_ulogic;
    OBDIV4       : in    std_ulogic;
    OBMUX0       : in    std_ulogic;
    OBMUX1       : in    std_ulogic;
    OBMUX2       : in    std_ulogic;
    DLYYB0       : in    std_ulogic;
    DLYYB1       : in    std_ulogic;
    DLYYB2       : in    std_ulogic;
    DLYYB3       : in    std_ulogic;
    DLYYB4       : in    std_ulogic;
    DLYGLB0      : in    std_ulogic;
    DLYGLB1      : in    std_ulogic;
    DLYGLB2      : in    std_ulogic;
    DLYGLB3      : in    std_ulogic;
    DLYGLB4      : in    std_ulogic;
    OCDIV0       : in    std_ulogic;
    OCDIV1       : in    std_ulogic;
    OCDIV2       : in    std_ulogic;
    OCDIV3       : in    std_ulogic;
    OCDIV4       : in    std_ulogic;
    OCMUX0       : in    std_ulogic;
    OCMUX1       : in    std_ulogic;
    OCMUX2       : in    std_ulogic;
    DLYYC0       : in    std_ulogic;
    DLYYC1       : in    std_ulogic;
    DLYYC2       : in    std_ulogic;
    DLYYC3       : in    std_ulogic;
    DLYYC4       : in    std_ulogic;
    DLYGLC0      : in    std_ulogic;
    DLYGLC1      : in    std_ulogic;
    DLYGLC2      : in    std_ulogic;
    DLYGLC3      : in    std_ulogic;
    DLYGLC4      : in    std_ulogic;
    FINDIV0      : in    std_ulogic;
    FINDIV1      : in    std_ulogic;
    FINDIV2      : in    std_ulogic;
    FINDIV3      : in    std_ulogic;
    FINDIV4      : in    std_ulogic;
    FINDIV5      : in    std_ulogic;
    FINDIV6      : in    std_ulogic;
    FBDIV0       : in    std_ulogic;
    FBDIV1       : in    std_ulogic;
    FBDIV2       : in    std_ulogic;
    FBDIV3       : in    std_ulogic;
    FBDIV4       : in    std_ulogic;
    FBDIV5       : in    std_ulogic;
    FBDIV6       : in    std_ulogic;
    FBDLY0       : in    std_ulogic;
    FBDLY1       : in    std_ulogic;
    FBDLY2       : in    std_ulogic;
    FBDLY3       : in    std_ulogic;
    FBDLY4       : in    std_ulogic;
    FBSEL0       : in    std_ulogic;
    FBSEL1       : in    std_ulogic;
    XDLYSEL      : in    std_ulogic;
    VCOSEL0      : in    std_ulogic;
    VCOSEL1      : in    std_ulogic;
    VCOSEL2      : in    std_ulogic;
    GLAOUT       : out   std_ulogic;
    LOCKOUT      : out   std_ulogic;
    GLBOUT       : out   std_ulogic;
    YBOUT        : out   std_ulogic;
    GLCOUT       : out   std_ulogic;
    YCOUT        : out   std_ulogic;
    VCOOUT       : out   std_ulogic
   );

  attribute VITAL_LEVEL0 of PLL_SDF : entity is TRUE;
end PLL_SDF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of PLL_SDF is
attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

constant PLL_pw_param : time := 1000.0/( VCOFREQUENCY * 2.0) * 1 ns;

signal CLKA_ipd               : std_ulogic;
  signal EXTFB_ipd              : std_ulogic;
  signal INTFB_ipd              : std_ulogic;
  signal POWERDOWN_ipd          : std_ulogic;

  signal AOUT                   : std_logic := 'X';
  signal BOUT                   : std_logic := 'X';
  signal COUT                   : std_logic := 'X';

  signal PLLCLK                 : std_logic := 'X';      -- PLL Core Output Clock 
                                                         -- with DIVN and DIVM applied
  signal CLKA_period            : Time      := 0.000 ns; -- Current CLKA period
  signal INTFB_period            : Time      := 0.000 ns; -- Current INTFB period

  signal PLLCLK_pw              : Time      := 10.0 ns; -- PLLCLK pulse width
  signal PLLCLK_period          : Time      := 10.0 ns;

  signal DIVN                   : Integer := 1; -- Divide by N divisor - range 1 to 128
  signal DIVM                   : Integer := 1; -- Multiply by M multiplier - range 1 to 128
  signal DIVU                   : Integer := 1; -- Divide by U divisor - range 1 to 32
  signal DIVV                   : Integer := 1; -- Divide by V divisor - range 1 to 32
  signal DIVW                   : Integer := 1; -- Divide by W divisor - range 1 to 32
  signal fb_loop_div            : Integer := 1; -- Total division of feedback loop

  signal CLKA2X                 : std_logic := 'X';

  signal UIN                    : std_logic := 'X'; -- Output of MUXA
  signal VIN                    : std_logic := 'X'; -- Output of MUXB
  signal WIN                    : std_logic := 'X'; -- Output of MUXC

  signal FBSEL                  : std_logic_vector( 1 downto 0 ) := "XX";
  signal FBSEL_illegal          : Boolean := False; -- True when FBSEL = 00

  signal OAMUX_config           : integer := -1;
  signal OBMUX_config           : integer := -1;
  signal OCMUX_config           : integer := -1;

  signal internal_lock          : boolean   := false;
  signal fin_period             : Time      := 0.000 ns;
  signal extfbin_fin_drift      : time      := 0 ps;
  signal locked                 : std_logic := '0'; -- 1 when PLL is externally locked as well as internally locked
  signal dly_locked                 : std_logic := '0';
  signal locked_vco0_edges      : integer   := -1;
  signal vco0_divu              : std_logic := '0';
  signal vco0_divv              : std_logic := '0';
  signal vco0_divw              : std_logic := '0';
  signal fin                    : std_logic := '0';
  signal CLKA_period_stable     : boolean   := false;
  signal INTFB_period_stable     : boolean   := false;
  signal EXTFB_period_stable     : boolean   := false;
  signal using_EXTFB            : std_logic := 'X';
  signal using_INTFB            : std_logic := 'X';
  signal EXTFB_delay_dtrmd      : Boolean   := false;
  signal calibrate_EXTFB_delay  : std_logic := '0';
  signal GLA_free_running       : std_logic := '1';
  signal AOUT_using_EXTFB       : std_logic := '1';
  signal GLA_pw                 : time      := 10.0 ns; -- Only used for external feedback
  signal EXTFB_period           : time      := 20.0 ns;  -- Only meaningful for external feedback
  signal external_dly_correct   : std_logic := 'X';

  signal internal_fb_delay      : time      := 0.000 ns;
  signal external_fb_delay      : time      := 0.000 ns;
  signal fb_delay      : time      := 0.000 ns;
  signal EXTFB_dly_dtrmd      : Boolean   := false;
  signal INTFB_dly_dtrmd      : Boolean   := false;
  signal fb_dly_dtrmd      : Boolean   := false;
signal vcoout_int            : std_logic := 'X';
signal final_lock            : std_logic;


  -- Use this instead of CONV_INTEGER to avoid ambiguous warnings
  function ulogic2int(
    vec  : std_ulogic_vector )
    return integer is
    variable result : integer;
    variable i : integer;
  begin
    result := 0;
    for i in vec'range loop
      result := result * 2;
      if vec(i) = '1' then
        result := result + 1;
      end if;
    end loop;
    return result;
  end function ulogic2int;

  function output_mux_driver( 
    outmux      : integer;
    halved      : std_logic;
    bypass      : std_logic;
    bypass2x    : std_logic;
    vco         : std_logic )
    return std_logic is
    variable result : std_logic;
  begin
     case outmux is
        when 1  => if ( '1' = halved ) then
                          result := bypass2x;
                       elsif ( '0' = halved ) then
                          result := bypass;
                       else
                          result := 'X';
                       end if;
        when 2  => result := vco;
        when 4  => result := vco;
        when 5  => result := vco;
        when 6  => result := vco;
        when 7  => result := vco;
        when others => result := 'X';
     end case;
     return result;
  end function output_mux_driver;

  begin

    ---------------------
    --  INPUT PATH DELAYs
    ---------------------
    WireDelay : block

    begin

      VitalWireDelay ( CLKA_ipd,      CLKA,      tipd_CLKA      );
      VitalWireDelay ( EXTFB_ipd,     EXTFB,     tipd_EXTFB     );
      VitalWireDelay ( INTFB_ipd,     INTFB,     tipd_INTFB     );
      VitalWireDelay ( POWERDOWN_ipd, POWERDOWN, tipd_POWERDOWN );
 
    end block WireDelay;

    -- #########################################################
    -- # Behavior Section
    -- #########################################################

    OAMUX_config <= ulogic2int( OAMUX2 & OAMUX1 & OAMUX0 );
    OBMUX_config <= ulogic2int( OBMUX2 & OBMUX1 & OBMUX0 );
    OCMUX_config <= ulogic2int( OCMUX2 & OCMUX1 & OCMUX0 );
    FBSEL <= TO_X01( FBSEL1 & FBSEL0 );

          LOCKOUT <= final_lock;

    DIVM <= ulogic2int( FBDIV6 & FBDIV5 & FBDIV4 & FBDIV3 & 
                        FBDIV2 & FBDIV1 & FBDIV0 ) + 1;

    DIVN <= ulogic2int( FINDIV6 & FINDIV5 & FINDIV4 & FINDIV3 & 
                        FINDIV2 & FINDIV1 & FINDIV0 ) + 1;

    DIVU <= ulogic2int( OADIV4 & OADIV3 & OADIV2 & OADIV1 & OADIV0 ) + 1;

    DIVV <= ulogic2int( OBDIV4 & OBDIV3 & OBDIV2 & OBDIV1 & OBDIV0 ) + 1;

    DIVW <= ulogic2int( OCDIV4 & OCDIV3 & OCDIV2 & OCDIV1 & OCDIV0 ) + 1;

    check_FBSEL : process
    begin
      wait on FBSEL, OAMUX_config, OBMUX_config, OCMUX_config, DIVM, DIVU, DIVN, CLKA_period_stable, PLLCLK_period, external_fb_delay;
      if ( IS_X( FBSEL ) ) then
         FBSEL_illegal <= true;
         assert ( not FBSEL'event )
            report "Warning: FBSEL is unknown." 
            severity Warning;
      elsif ( "00" = FBSEL ) then -- Grounded.
         FBSEL_illegal <= true;
         assert ( not FBSEL'event )
            report "Warning: Illegal FBSEL configuration 00." 
            severity Warning;
      elsif ( "11" = FBSEL ) then -- External feedback
         if ( 2 > OAMUX_config ) then
            FBSEL_illegal <= true;
            assert  ( not ( FBSEL'event or OAMUX_config'event ) )
               report "Illegal configuration. GLA cannot be in bypass mode (OAMUX = 000 or OAMUX = 001) when using external feedback (FBSEL = 11)." 
               severity Warning;
         elsif ( DIVM < 5 ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or DIVM'event ) )
               report "Error: FBDIV must be greater than 4 when using external feedback (FBSEL = 11)."
               severity Error;
         elsif ( ( DIVM * DIVU ) > 232 ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or DIVM'event or DIVU'event ) )
               report "Error: Product of FBDIV and OADIV must be less than 233 when using external feedback (FBSEL = 11)."
               severity Error;
         elsif ( ( DIVN mod DIVU ) /= 0 ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or DIVN'event or DIVU'event ) )
               report "Error: Division factor FINDIV must be a multiple of OADIV when using external feedback (FBSEL = 11)."
               severity Error;
         elsif ( CLKA_period_stable and EXTFB_delay_dtrmd and
                 ( ( 1 < OBMUX_config ) or ( 1 < OCMUX_config ) ) and
                 ( ( external_fb_delay >= CLKA_period ) or ( external_fb_delay >= PLLCLK_period ) ) ) then
            FBSEL_illegal <= true;
            assert ( not ( FBSEL'event or CLKA_period_stable'event or external_fb_delay'event or PLLCLK_period'event ) )
              report "Error: Total sum of delays in the feedback path must be less than 1 VCO period AND less than 1 CLKA period when V and/or W dividers when using external feedback (FBSEL = 11)."
               severity Error;
         else
            FBSEL_illegal <= false;
         end if;
      else
         FBSEL_illegal <= false;
      end if;
    end process check_FBSEL;

    -- Mimicing silicon - no need for a 50/50 duty cycle and this way fin only changes on rising edge of CLKA (except when DIVN is 1)
    gen_fin: process
      variable num_CLKA_re   : integer;
    begin
       wait until rising_edge( CLKA_ipd );
       fin <= '1';
       num_CLKA_re := 0;
       while ( 'X' /= TO_X01( CLKA_ipd ) ) loop
          wait on CLKA_ipd;
          if ( 1 = DIVN )then
             fin <= CLKA_ipd;
          elsif ( '1' = CLKA_ipd ) then
             num_CLKA_re := num_CLKA_re + 1;
             if ( ( num_CLKA_re mod DIVN  ) = 0 ) then
                fin <= '1';
                num_CLKA_re := 0;
             elsif ( ( num_CLKA_re mod DIVN ) = 1 ) then
                fin <= '0';
             end if;
          end if;
       end loop;
    end process gen_fin;

--    PLL_pw_param <=  1000.0/real(VCOFREQUENCY) * 1 ns;
    
    gen_vcoout: process
      begin
        vcoout_int <= '1';
        wait for PLL_pw_param;
        vcoout_int <= '0';
        wait for PLL_pw_param;        
      end process gen_vcoout;

      VCOOUT <= vcoout_int;
      
    GetINTFBPeriod : process ( INTFB_ipd, POWERDOWN_ipd )
      variable re                 : Time :=  0.000 ns; -- Current INTFB rising edge
      variable INTFB_num_re_stable : Integer := -1;  
    begin
      if ( TO_X01( POWERDOWN_ipd ) = '1' )  then
        if ( INTFB_ipd'event and ( '1' = TO_X01( INTFB_ipd ) ) ) then
           if ( INTFB_period /= ( NOW - re ) ) then
              INTFB_period <= ( NOW - re );
              INTFB_num_re_stable := -1;
              INTFB_period_stable <= false;
           else
             if ( 3 > INTFB_num_re_stable ) then
               INTFB_num_re_stable := INTFB_num_re_stable + 1;
             elsif ( 3 = INTFB_num_re_stable ) then
               INTFB_period_stable <= true;
             end if;
           end if;
           re := NOW;
        elsif ( INTFB_period < ( NOW - re ) ) then
           INTFB_num_re_stable := -1;
           INTFB_period_stable <= false;
        end if;
      else
        INTFB_num_re_stable := -1;
        INTFB_period_stable <= false;
      end if;
    end process GetINTFBPeriod;

    calc_internal_fb_delay : process
      variable vco_re : time;
      variable internal_fb_re : time;
      variable tmp_internal_delay : time;
    begin
      intfb_dly_dtrmd <= false;
      wait until (INTFB_period_stable = true );      
      wait until rising_edge( vcoout_int );
      wait until rising_edge( vcoout_int );
      vco_re := NOW;        
      wait until rising_edge( INTFB_ipd );
      internal_fb_re := NOW;
      tmp_internal_delay := internal_fb_re - vco_re;
      if (tmp_internal_delay = INTFB_period) then
        tmp_internal_delay := 0 ns;
      end if;
      internal_fb_delay <= tmp_internal_delay;
      intfb_dly_dtrmd <= true;
      wait until INTFB_period_stable = false;
    end process calc_internal_fb_delay;

   GetEXTFBPeriod : process ( EXTFB_ipd, POWERDOWN_ipd )
      variable re                 : Time :=  0.000 ns; -- Current EXTFB rising edge
      variable EXTFB_num_re_stable : Integer := -1;  
    begin
      if ( TO_X01( POWERDOWN_ipd ) = '1' )  then
        if ( EXTFB_ipd'event and ( '1' = TO_X01( EXTFB_ipd ) ) ) then
           if ( EXTFB_period /= ( NOW - re ) ) then
              EXTFB_period <= ( NOW - re );
              EXTFB_num_re_stable := -1;
              EXTFB_period_stable <= false;
           else
             if ( 3 > EXTFB_num_re_stable ) then
               EXTFB_num_re_stable := EXTFB_num_re_stable + 1;
             elsif ( 3 = EXTFB_num_re_stable ) then
               EXTFB_period_stable <= true;
             end if ;
           end if;
           re := NOW;
        elsif ( EXTFB_period < ( NOW - re ) ) then
           EXTFB_num_re_stable := -1;
           EXTFB_period_stable <= false;
        end if;
      else
        EXTFB_num_re_stable := -1;
        EXTFB_period_stable <= false;
      end if;
    end process GetEXTFBPeriod;

     calc_external_fb_delay : process 
      variable clka_fb_re : time := 0.000 ns;
      variable external_fb_re : time := 0.000 ns;
      variable tmp_external_delay : time := 0.000 ns;
    begin
      extfb_dly_dtrmd <= false;
      wait until (using_EXTFB = '1' and CLKA_period_stable = true);
      wait until rising_edge( CLKA_ipd );
      clka_fb_re := NOW;        
      wait until rising_edge( EXTFB_ipd );
      external_fb_re := NOW;
      tmp_external_delay := external_fb_re - clka_fb_re;
      if (tmp_external_delay = INTFB_period or
          tmp_external_delay = CLKA_period) then
        tmp_external_delay := 0 ns;
      end if;
      external_fb_delay <= tmp_external_delay;
      extfb_dly_dtrmd <= true;
      wait until falling_edge (dly_locked);
    end process calc_external_fb_delay;     

      select_fb_delay: process (external_fb_delay, internal_fb_delay)
      begin  -- process select_fb_delay
        if (using_EXTFB = '1') then
          fb_delay <= external_fb_delay;
        else
          fb_delay <= internal_fb_delay;          
        end if;  
      end process select_fb_delay;

      fb_dly_dtrmd <= extfb_dly_dtrmd when using_EXTFB = '1'
                      else intfb_dly_dtrmd;
        
    GetCLKAPeriod : process ( CLKA_ipd, POWERDOWN_ipd, FBSEL_illegal, locked_vco0_edges, external_dly_correct )
      -- locked_vco0_edges is in the sensitivity list so that we periodically check for CLKA stopped
      variable re                 : Time :=  0.000 ns; -- Current CLKA rising edge
      variable CLKA_num_re_stable : Integer := -1;   -- Number of CLKA rising edges that PLL config stable
    begin
      if (( TO_X01( POWERDOWN_ipd ) = '1' ) and ( FBSEL_illegal = False ))  then
        if ( CLKA_ipd'event and ( '1' = TO_X01( CLKA_ipd ) ) ) then
           if ( CLKA_period /= ( NOW - re ) ) then
              CLKA_period <= ( NOW - re );
              CLKA_num_re_stable := -1;
              internal_lock <= false;
              CLKA_period_stable <= false;
           else
              if ( f_CLKA_LOCK > CLKA_num_re_stable ) then
                 CLKA_num_re_stable := CLKA_num_re_stable + 1;
              elsif ( f_CLKA_LOCK = CLKA_num_re_stable and fb_dly_dtrmd = true) then
                 internal_lock <=  true;
              end if;
              CLKA_period_stable <= true;
           end if;
           re := NOW;
        elsif ( CLKA_period < ( NOW - re ) ) then
           CLKA_num_re_stable := -1;
           internal_lock <= false;
           CLKA_period_stable <= false;
        end if;
      else
        CLKA_num_re_stable := -1;
        internal_lock <= false;
        CLKA_period_stable <= false;
      end if;
    end process GetCLKAPeriod;

    fin_period         <= CLKA_period * DIVN;

    GLA_pw             <= PLLCLK_pw * DIVU;

    extfbin_fin_drift  <= ( GLA_pw * DIVM * 2.0 ) - fin_period;

    PLLCLK_period      <= fin_period / real( fb_loop_div );

    PLLCLK_pw          <= PLLCLK_period / 2.0;

    calc_fb_loop_div : process( DIVM, DIVU, using_EXTFB )
    begin
       if ( using_EXTFB  = '1' ) then
           fb_loop_div <= DIVM * DIVU; 
       else
           fb_loop_div <= DIVM;
       end if;
    end process calc_fb_loop_div;

    sync_pll : process( fin, internal_lock )
    begin
       if ( not( internal_lock ) ) then
          locked <= '0';
       elsif ( rising_edge( fin ) ) then
          locked <= '1';
       end if;
    end process sync_pll;

     dly_locked <= transport locked after ( CLKA_period - fb_delay );

      gen_lock : process( CLKA_ipd, POWERDOWN_ipd)
        begin
          if ( TO_X01(POWERDOWN_ipd) = '0') then
            final_lock <= '0';
            elsif ( TO_X01(CLKA_ipd) = 'X' ) then
              final_lock <= 'X';
            elsif rising_edge (CLKA_ipd) then                            
                final_lock <= locked;
          end if;
        end process gen_lock;
        
    count_locked_vco0_edges: process( dly_locked, locked_vco0_edges )
    begin
       if ( dly_locked'event ) then
          if ( dly_locked = '1' ) then
            locked_vco0_edges <= 0;
          else
            locked_vco0_edges <= -1;
          end if;
       elsif ( dly_locked = '1' ) then
          if ( ( locked_vco0_edges mod( DIVU * DIVV * DIVW * DIVM * 2 ) ) = 0 ) then
             locked_vco0_edges <= 1 after PLLCLK_pw;
          else
             locked_vco0_edges <= ( locked_vco0_edges + 1 ) after PLLCLK_pw;
          end if;
       end if;
    end process count_locked_vco0_edges;

    gen_vco0_div: process( locked_vco0_edges )
    begin
       if ( locked_vco0_edges = -1 ) then
          vco0_divu <= '0';
          vco0_divv <= '0';
          vco0_divw <= '0';
       else 
         if ( ( locked_vco0_edges mod DIVU ) = 0 ) then
           vco0_divu <= not vco0_divu;
         end if;
         if ( ( locked_vco0_edges mod DIVV ) = 0 ) then
           vco0_divv <= not vco0_divv;
         end if;
         if ( ( locked_vco0_edges mod DIVW ) = 0 ) then
           vco0_divw <= not vco0_divw;
         end if;
       end if;
    end process gen_vco0_div;

    UIN <= output_mux_driver(  OAMUX_config, '0', CLKA_ipd, CLKA2X, vco0_divu );
    VIN <= output_mux_driver(  OBMUX_config, '0', '0', '0', vco0_divv );
    WIN <= output_mux_driver(  OCMUX_config, '0', '0', '0', vco0_divw );

    double_CLKA: process( CLKA_ipd )
       variable re      : Time := 0 ns;
       variable prev_re : Time := 0 ns;
       variable period  : Time := 0 ns;
    begin
       if ( TO_X01( CLKA_ipd ) = '1' ) then
         prev_re := re;
         re := NOW;
         period := re - prev_re;
         if ( period > 0 ns ) then
            CLKA2X <= '1';
            CLKA2X <= transport '0' after ( period / 4.0 );
            CLKA2X <= transport '1' after ( period / 2.0 );
            CLKA2X <= transport '0' after ( period * 3.0 / 4.0 );
         end if;
       end if;
    end process double_CLKA;

    --
    -- AOUT Output of Divider U
    --

    DividerU : process ( UIN, CLKA_ipd, POWERDOWN_ipd )

      variable force_0         : Boolean  := True;
      variable num_edges       : Integer  := -1;
      variable res_post_reset1 : Integer  :=  0;
      variable fes_post_reset1 : Integer  :=  0;
      variable res_post_reset0 : Integer  :=  0;
      variable fes_post_reset0 : Integer  :=  0;

    begin

      if ( 1 = OAMUX_config ) then -- PLL core bypassed.  OADIVRST active.

        if ( CLKA_ipd'event ) then
          if ( TO_X01( CLKA_ipd ) = '1' and TO_X01( CLKA_ipd'last_value ) = '0' ) then
             if ( 4 > res_post_reset1 ) then
                res_post_reset1 := res_post_reset1 + 1;
             end if;
             if ( 4 > res_post_reset0 ) then
               res_post_reset0 := res_post_reset0 + 1;
             end if;
             if ( res_post_reset1 = 3 ) then
                force_0 := False;
                num_edges := -1;
             end if;
          elsif ( TO_X01( CLKA_ipd ) = '0' and TO_X01( CLKA_ipd'last_value ) = '1' ) then
             if ( 4 > fes_post_reset1 ) then
               fes_post_reset1 := fes_post_reset1 + 1;
             end if;
             if ( 4 > fes_post_reset0 ) then
               fes_post_reset0 := fes_post_reset0 + 1;
             end if;
             if ( fes_post_reset1 = 1 ) then
                force_0 := True;
             end if;
          end if;
        end if;

        if ( UIN'event ) then
          num_edges := num_edges + 1;
          if ( force_0 ) then
            AOUT <= '0';
          elsif ( TO_X01( UIN ) = 'X' ) then
            AOUT <= 'X';
          elsif ( ( num_edges mod DIVU ) = 0 ) then
            num_edges := 0;
            if ( TO_X01 ( AOUT ) = 'X' ) then
              AOUT <= UIN;
            else
              AOUT <= not AOUT;
            end if;
          end if;
        end if;

      else -- PLL not bypassed
        if ( TO_X01 ( POWERDOWN_ipd ) = '0' ) then
          AOUT <= '0';
        elsif ( TO_X01 ( POWERDOWN_ipd ) = '1' ) then
          AOUT <= UIN;
        else -- POWERDOWN unknown
          AOUT <= 'X';
        end if;
      end if;

    end process DividerU;


    --
    -- BOUT Output of Divider V
    --

    DividerV : process ( VIN, POWERDOWN_ipd )

      variable force_0         : Boolean  := True;
      variable num_edges       : Integer  := -1;
      variable res_post_reset1 : Integer  :=  0;
      variable fes_post_reset1 : Integer  :=  0;
      variable res_post_reset0 : Integer  :=  0;
      variable fes_post_reset0 : Integer  :=  0;

    begin

      if ( 0 = OBMUX_config ) then
        BOUT <= 'X';
      elsif ( 1 = OBMUX_config ) then -- PLL core bypassed.  OBDIVRST active.
        if ( VIN'event ) then
          num_edges := num_edges + 1;
          if ( force_0 ) then
            BOUT <= '0';
          elsif ( TO_X01( VIN ) = 'X' ) then
            BOUT <= 'X';
          elsif ( ( num_edges mod DIVV ) = 0 ) then
            num_edges := 0;
            if ( TO_X01 ( BOUT ) = 'X' ) then
              BOUT <= VIN;
            else
              BOUT <= not BOUT;
            end if;
          end if;
        end if;
      else -- PLL not bypassed
        if ( TO_X01 ( POWERDOWN_ipd ) = '0' ) then
          BOUT <= '0';
        elsif ( TO_X01 ( POWERDOWN_ipd ) = '1' ) then
          BOUT <= VIN;
        else -- POWERDOWN unknown
          BOUT <= 'X';
        end if;
      end if;

    end process DividerV;

    --
    -- COUT Output of Divider W
    --

    DividerW : process ( WIN, POWERDOWN_ipd )

      variable force_0         : Boolean  := True;
      variable num_edges       : Integer  := -1;
      variable res_post_reset1 : Integer  :=  0;
      variable fes_post_reset1 : Integer  :=  0;
      variable res_post_reset0 : Integer  :=  0;
      variable fes_post_reset0 : Integer  :=  0;

    begin

      if ( 0 = OCMUX_config ) then
        COUT <= 'X';
      elsif ( 1 = OCMUX_config ) then -- PLL core bypassed.  OCDIVRST active.
        if ( WIN'event ) then
          num_edges := num_edges + 1;
          if ( force_0 ) then
            COUT <= '0';
          elsif ( TO_X01( WIN ) = 'X' ) then
            COUT <= 'X';
          elsif ( ( num_edges mod DIVW ) = 0 ) then
            num_edges := 0;
            if ( TO_X01 ( COUT ) = 'X' ) then
              COUT <= WIN;
            else
              COUT <= not COUT;
            end if;
          end if;
        end if;

      else -- PLL not bypassed
        if ( TO_X01 ( POWERDOWN_ipd ) = '0' ) then
          COUT <= '0';
        elsif ( TO_X01 ( POWERDOWN_ipd ) = '1' ) then
          COUT <= WIN;
        else -- POWERDOWN unknown
          COUT <= 'X';
        end if;
      end if;

    end process DividerW;

    using_EXTFB <= TO_X01( FBSEL1 and FBSEL0 );

--    external_dly_correct <= expected_EXTFB xnor EXTFB_ipd after 1 ps;

    Aoutputs: process( AOUT, CLKA_ipd, OAMUX_config  )
    begin
        if ( 0 = OAMUX_config ) then
          GLAOUT <=  CLKA_ipd;
        elsif ( ( 1 = OAMUX_config ) or ( 3 = OAMUX_config ) ) then
          GLAOUT <= 'X';
          assert ( not OAMUX_config'event )
            report "WARNING: Illegal OAMUX configuration."
            severity warning; 
        elsif (fb_dly_dtrmd = false and using_EXTFB = '1') then
          GLAOUT <= CLKA_ipd;
        else                                              
          GLAOUT <= AOUT;
        end if;
    end process Aoutputs;
    
    Boutputs: process ( BOUT, OBMUX_config )
    begin
      if ( ( 0 = OBMUX_config ) or ( 1 = OBMUX_config ) or
           ( 3 = OBMUX_config ) ) then
          GLBOUT <=  'X';
          YBOUT  <=  'X';
          assert ( not OBMUX_config'event )
            report "WARNING: Illegal OBMUX configuration."
            severity warning;
        else
          GLBOUT <=  BOUT;
          YBOUT  <=  BOUT;
        end if;
    end process Boutputs;

    Coutputs: process ( COUT, OCMUX_config )
    begin
      if ( ( 0 = OCMUX_config ) or ( 1 = OCMUX_config ) or
           ( 3 = OCMUX_config ) ) then
        GLCOUT <=  'X';
        YCOUT  <=  'X';
          assert ( not OCMUX_config'event )
            report "WARNING: Illegal OCMUX configuration."
            severity warning;
        else
          GLCOUT <=  COUT;
          YCOUT  <=  COUT;
        end if;
    end process Coutputs;
    
  end VITAL_ACT;

configuration CFG_PLL_SDF_VITAL of PLL_SDF is
  for VITAL_ACT
  end for;
end CFG_PLL_SDF_VITAL;
--***************************************************************************
--***************************************************************************
-- Detailed Revision History:
--
-- Version  Date(MM/DD/YY)   Submitter              Description
--
-- 1.0      10/8/09         Kiran Yerribandi     First Version.
--------------------------------------------------------------------
--------------------------------------------------------------------
-- CELL NAME : PLL_DLY_SDF
---------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity PLL_DLY_SDF is
  generic (
    VCOFREQUENCY       :  Real    := 0.0;
    InstancePath       :  String           := "*";
    Xon                :  Boolean          := False;
    MsgOn              :  Boolean          := True;
    tpd_GLAIN_GLA          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_GLBIN_GLB          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_GLCIN_GLC          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_YBIN_YB          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_YCIN_YC          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_LOCKIN_LOCK          :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_EXTFBIN_EXTFBOUT         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns );
    tpd_VCOIN_PLLOUT         :  VitalDelayType01 := ( 0.000 ns, 0.000 ns )
    );
  port (
    GLAIN  : in  std_ulogic;
    GLBIN  : in  std_ulogic;
    GLCIN  : in  std_ulogic;
    YBIN  : in  std_ulogic;
    YCIN  : in  std_ulogic;
    VCOIN  : in  std_ulogic;
    LOCKIN  : in  std_ulogic;
    EXTFBIN  : in  std_ulogic;
    GLA : out std_ulogic;
    GLB : out std_ulogic;
    GLC : out std_ulogic;
    YB : out std_ulogic;
    YC : out std_ulogic;
    PLLOUT : out std_ulogic;
    LOCK : out std_ulogic;    
    EXTFBOUT : out std_ulogic);

  attribute VITAL_LEVEL0 of PLL_DLY_SDF : entity is TRUE;
end PLL_DLY_SDF;

library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of PLL_DLY_SDF is
  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;
begin

  gla_process : process (GLAIN)
    variable GLA_zd : std_ulogic;
    variable GLA_GlitchData : VitalGlitchDataType;
  begin

    GLA_zd := TO_X01(GLAIN);

    VitalPathDelay01 (
      OutSignal => GLA,
      GlitchData => GLA_GlitchData,
      OutSignalName => "GLA",
      OutTemp => GLA_zd,
      Paths => (
        0 => (GLAIN'last_event,tpd_GLAIN_GLA, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;


  glb_process : process (GLBIN)
    variable GLB_zd : std_ulogic;
    variable GLB_GlitchData : VitalGlitchDataType;
  begin

    GLB_zd := TO_X01(GLBIN);

    VitalPathDelay01 (
      OutSignal => GLB,
      GlitchData => GLB_GlitchData,
      OutSignalName => "GLB",
      OutTemp => GLB_zd,
      Paths => (
        0 => (GLBIN'last_event,tpd_GLBIN_GLB, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;


  glc_process : process (GLCIN)
    variable GLC_zd : std_ulogic;
    variable GLC_GlitchData : VitalGlitchDataType;
  begin

    GLC_zd := TO_X01(GLCIN);

    VitalPathDelay01 (
      OutSignal => GLC,
      GlitchData => GLC_GlitchData,
      OutSignalName => "GLC",
      OutTemp => GLC_zd,
      Paths => (
        0 => (GLCIN'last_event,tpd_GLCIN_GLC, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;


  yb_process : process (YBIN)
    variable YB_zd : std_ulogic;
    variable YB_GlitchData : VitalGlitchDataType;
  begin

    YB_zd := TO_X01(YBIN);

    VitalPathDelay01 (
      OutSignal => YB,
      GlitchData => YB_GlitchData,
      OutSignalName => "YB",
      OutTemp => YB_zd,
      Paths => (
        0 => (YBIN'last_event,tpd_YBIN_YB, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;


  yc_process : process (YCIN)
    variable YC_zd : std_ulogic;
    variable YC_GlitchData : VitalGlitchDataType;
  begin

    YC_zd := TO_X01(YCIN);

    VitalPathDelay01 (
      OutSignal => YC,
      GlitchData => YC_GlitchData,
      OutSignalName => "YC",
      OutTemp => YC_zd,
      Paths => (
        0 => (YCIN'last_event,tpd_YCIN_YC, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;


  lock_process : process (LOCKIN)
    variable LOCK_zd : std_ulogic;
    variable LOCK_GlitchData : VitalGlitchDataType;
  begin

    LOCK_zd := TO_X01(LOCKIN);

    VitalPathDelay01 (
      OutSignal => LOCK,
      GlitchData => LOCK_GlitchData,
      OutSignalName => "LOCK",
      OutTemp => LOCK_zd,
      Paths => (
        0 => (LOCKIN'last_event,tpd_LOCKIN_LOCK, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;


  vco_process : process (VCOIN)
    variable PLLOUT_zd : std_ulogic;
    variable PLLOUT_GlitchData : VitalGlitchDataType;
  begin

    PLLOUT_zd := TO_X01(VCOIN);

    VitalPathDelay01 (
      OutSignal => PLLOUT,
      GlitchData => PLLOUT_GlitchData,
      OutSignalName => "PLLOUT",
      OutTemp => PLLOUT_zd,
      Paths => (
        0 => (VCOIN'last_event,tpd_VCOIN_PLLOUT, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;

 
  extfb_process : process (EXTFBIN)
    variable EXTFBOUT_zd : std_ulogic;
    variable EXTFBOUT_GlitchData : VitalGlitchDataType;
  begin

    EXTFBOUT_zd := TO_X01(EXTFBIN);

    VitalPathDelay01 (
      OutSignal => EXTFBOUT,
      GlitchData => EXTFBOUT_GlitchData,
      OutSignalName => "EXTFBOUT",
      OutTemp => EXTFBOUT_zd,
      Paths => (
        0 => (EXTFBIN'last_event,tpd_EXTFBIN_EXTFBOUT, true)),
      Mode => VitalTransport,
      Xon => Xon,
      MsgOn => MsgOn,
      MsgSeverity => WARNING);    
    
  end process;
  
end VITAL_ACT;

configuration CFG_PLL_DLY_SDF_VITAL of PLL_DLY_SDF is
  for VITAL_ACT
  end for;
end CFG_PLL_DLY_SDF_VITAL;
