-- -------------------------------------------------------------------- 
-- >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<< 
-- -------------------------------------------------------------------- 
-- Copyright (c) 2005 by Lattice Semiconductor Corporation 
-- -------------------------------------------------------------------- 
-- 
-- 
--                     Lattice Semiconductor Corporation 
--                     5555 NE Moore Court 
--                     Hillsboro, OR 97214 
--                     U.S.A 
-- 
--                     TEL: 1-800-Lattice (USA and Canada) 
--                          408-826-6000 (other locations) 
-- 
--                     web: http://www.latticesemi.com/ 
--                     email: techsupport@latticesemi.com 
-- 
-- 
-- Revision History : 

--***************************************************************
--	This VHDL file contains the source code of the complete
--	library modules in a single file  including the lattice 
--	declaration package which contains the declaration and 
--  instantiation of the primitives
--***************************************************************

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE STD.TEXTIO.ALL;

package VHD_PKG is

	component SHFE 
		port( REF : IN std_logic;
			  DATA : IN std_logic);
	end component;

	component PW 
		port( PULSE : IN std_logic);
	end component;

	component INV 
		port( A0 : IN std_logic;
			  ZN0 : OUT std_logic);
	end component;

	component BUF 
		port( A0 : IN std_logic;
			  Z0 : OUT std_logic);
	end component;

	component LXOR2
		port(A0 : IN std_logic;
			 A1 : IN std_logic;
			 Z0 : OUT std_logic);
	end component;

	component FD11
		port(D0 : IN std_logic;
			 CLK : IN std_logic;
			 Q0 : OUT std_logic);
	end component;

	component FD21
		port(D0 : IN std_logic;
			 CLK : IN std_logic;
			 CD : IN std_logic;
			 Q0 : OUT std_logic);
	end component;

	component XINV 
		port( A0 : IN std_logic;
			  ZN0 : OUT std_logic);
	end component;

	component XINPUT 
		port( XI0 : IN std_logic;
			  Z0 : OUT std_logic);
	end component;

	component XOUTPUT 
		port( A0 : IN std_logic;
			  XO0 : OUT std_logic);
	end component;

	component XBIDI1 
		port ( A0 : IN std_logic;
			   OE : IN std_logic;
			   Z0 : OUT std_logic;
			   XB0 : INOUT std_logic);
	 end component;

	component XTRI1 
		port( A0 : IN  std_logic;
			  OE : IN  std_logic;
			  XO0 : OUT  std_logic);
	end component;

	component XDFF1
		port( D0 : IN std_logic;
			  CLK : IN std_logic;
			  Q0 : OUT std_logic);
	end component;

	component XDL1
		port ( D0 : IN std_logic;
				G : IN std_logic;
			   Q0 : OUT std_logic);
	end component;

component XOR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND13 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND14 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND15 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND17 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 A16 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND18 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 A16 : IN std_logic;
		 A17 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component NAND2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component FD11E
  port (D0, CLK, EN : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component FD21E
  port (D0, CLK, CD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component FDC1
  port (D0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component FDC1E
  port (D0, CLK, SD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component FDE1
  port (D0, CLK, CD, SD : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component FDE1E
  port (D0, CLK, CD, SD, EN : IN std_logic;
	               Q0 : OUT std_logic);
end component;

component FTI21
  port (T0, CLK, CD : IN std_logic;
                 Q0 : OUT std_logic);
end component;

component FTI21E
  port (T0, CLK, CD, EN : IN std_logic;
                     Q0 : OUT std_logic);
end component;

component FTI31
  port (T0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component FTI31E
  port (T0, CLK, SD, EN : IN std_logic;
		 Q0 : OUT std_logic);
end component;

component FTI41
  port (T0, CLK, SD, CD : IN std_logic;
		 Q0 : OUT std_logic);
end component;

component FTI41E
  port (T0, CLK, CD, SD, EN : IN std_logic;
		     Q0 : OUT std_logic);
end component;

component IT11
  port(A0, OE : IN std_logic;
	 O0 : OUT  std_logic);
end component;
       
component LDI11
  port (D0, G : IN std_logic;
           Q0 : OUT std_logic);
end component;

component LDI21
  port (D0, G, CD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component LDI31
  port (D0, G, SD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component LDI41
  port (D0, G, CD, SD : IN std_logic;
	         Q0 : OUT std_logic);
end component;

component XDFF1E
  port (D0, CLK, EN : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component XDFF2
  port (D0, CLK, CD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component XDFF2E
  port (D0, CLK, CD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component XDFF3
  port (D0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component XDFF3E
  port (D0, CLK, SD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component XDFF4
  port (D0, CLK, CD, SD : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component XDFF4E
  port (D0, CLK, CD, SD, EN : IN std_logic;
	               Q0 : OUT std_logic);
end component;

component XDL2
  port (D0, G, CD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component XDL3
  port (D0, G, SD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component XDL4
  port (D0, G, CD, SD : IN std_logic;
	         Q0 : OUT std_logic);
end component;

component ADDF1
  port (
    Z0 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic;
    CI : in std_logic);
end component;
component ADDF16A
  port (
    CO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic;
    CI : in std_logic);
end component;
component ADDF2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    CI : in std_logic);
end component;
component ADDF4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    CI : in std_logic);
end component;
component ADDF8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    CI : in std_logic);
end component;
component ADDF8A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    CI : in std_logic);
end component;
component ADDH1
  port (
    Z0 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic);
end component;
component ADDH16A
  port (
    CO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic);
end component;
component ADDH2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic);
end component;
component ADDH3
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic);
end component;
component ADDH4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component ADDH8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component ADDH8A
  port (
    CO : out std_logic;
    Z7 : out std_logic;
    Z6 : out std_logic;
    Z5 : out std_logic;
    Z4 : out std_logic;
    Z3 : out std_logic;
    Z2 : out std_logic;
    Z1 : out std_logic;
    Z0 : out std_logic;
    B7 : in std_logic;
    B6 : in std_logic;
    B5 : in std_logic;
    B4 : in std_logic;
    B3 : in std_logic;
    B2 : in std_logic;
    B1 : in std_logic;
    B0 : in std_logic;
    A7 : in std_logic;
    A6 : in std_logic;
    A5 : in std_logic;
    A4 : in std_logic;
    A3 : in std_logic;
    A2 : in std_logic;
    A1 : in std_logic;
    A0 : in std_logic);
end component;
component BI11
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI14
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI18
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BI21
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI28
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BI31
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI34
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI38
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BI41
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI48
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BIID11
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID11E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIID14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID14E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIID18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID21
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID31
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID41
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID51
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID61
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID71
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID81
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID91
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID91E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIID94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID94E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIIDA1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDA1E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDA4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB1E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIL11
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL21
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL31
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL41
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL51
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL61
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL71
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL81
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL91
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIILA1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIILA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIILB1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIILB4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIN27
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic);
end component;
component BIOD11
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component BIOD11E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD14
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component BIOD14E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD21
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component BIOD21E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component BIOD24E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD31
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD31E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD34
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD34E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD41
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD41E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD44E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL11
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL14
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL21
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL31
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL34
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL41
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component CBD11
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD12
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD21
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD22
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD31
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD32
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD41
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD42
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD516
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD616
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CAO : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD84
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBD88
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBD94
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBD98
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBDA16
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D10 : in std_logic;
    D11 : in std_logic;
    D12 : in std_logic;
    D13 : in std_logic;
    D14 : in std_logic;
    D15 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    D8 : in std_logic;
    D9 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDA4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDA8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDB4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDB8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBU11
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU12
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU21
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU22
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU31
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU32
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU41
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU42
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU516
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU616
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CAO : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU716
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D10 : in std_logic;
    D11 : in std_logic;
    D12 : in std_logic;
    D13 : in std_logic;
    D14 : in std_logic;
    D15 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    D8 : in std_logic;
    D9 : in std_logic;
    EN : in std_logic;
    LD : in std_logic);
end component;
component CBU84
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBU88
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBU94
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBU98
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBUA16
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D10 : in std_logic;
    D11 : in std_logic;
    D12 : in std_logic;
    D13 : in std_logic;
    D14 : in std_logic;
    D15 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    D8 : in std_logic;
    D9 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUA4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUA8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUB4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUB8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUD1
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD2
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD4S
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    DNUP : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUD8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD8S
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    DNUP : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CDD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDUD4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CDUD4C
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CDUD8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CDUD8C
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CGD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CGD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CGD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CGU14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CGU24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CGU34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CGUD4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CGUD4S
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    DNUP : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CMP2
  port (
    EQ : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic);
end component;
component CMP4
  port (
    EQ : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component CMP8
  port (
    EQ : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component DEC2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    S0 : in std_logic);
end component;
component DEC2E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DEC3
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DEC3E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DEC4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DEC4E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX22
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX22E
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DMUX24
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX24E
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX2E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DMUX4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX42
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX42E
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DMUX44
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    W2 : out std_logic;
    W3 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    X2 : out std_logic;
    X3 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX44E
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    W2 : out std_logic;
    W3 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    X2 : out std_logic;
    X3 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX4E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX82
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Y4 : out std_logic;
    Y5 : out std_logic;
    Y6 : out std_logic;
    Y7 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX82E
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Y4 : out std_logic;
    Y5 : out std_logic;
    Y6 : out std_logic;
    Y7 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component F3ADD
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    G012 : out std_logic;
    P012 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    CI : in std_logic);
end component;
component F3SUB
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    G012 : out std_logic;
    P012 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    BI : in std_logic);
end component;
component FD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic);
end component;
component FD14E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component FD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic);
end component;
component FD18E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic);
end component;
component FD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FD24E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component FD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FD28E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic);
end component;
component FD31
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic);
end component;
component FD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic);
end component;
component FD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic);
end component;
component FD41
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FD51
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component FD54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component FD58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component FD61
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FD64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FD68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FD71
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD81
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    TE : in std_logic);
end component;
component FD84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    TE : in std_logic);
end component;
component FD88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    TE : in std_logic);
end component;
component FD91
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD98
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FDA1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic;
    TE : in std_logic);
end component;
component FDA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic;
    TE : in std_logic);
end component;
component FDA8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic;
    TE : in std_logic);
end component;
component FDB1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    SD : in std_logic);
end component;
component FDB4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    SD : in std_logic);
end component;
component FDB8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    SD : in std_logic);
end component;
component FDC4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component FDC4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FDC8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    SD : in std_logic);
end component;
component FDC8E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FDE4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component FDE4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FDE8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    SD : in std_logic);
end component;
component FDE8E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FJK11
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    CLK : in std_logic);
end component;
component FJK21
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FJK31
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FJK41
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FJK51
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FJK61
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    SD : in std_logic);
end component;
component FJK64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    SD : in std_logic);
end component;
component FJK68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    J4 : in std_logic;
    J5 : in std_logic;
    J6 : in std_logic;
    J7 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    K4 : in std_logic;
    K5 : in std_logic;
    K6 : in std_logic;
    K7 : in std_logic;
    SD : in std_logic);
end component;
component FJK71
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    SD : in std_logic);
end component;
component FJK71E
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    SD : in std_logic);
end component;
component FJK74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    SD : in std_logic);
end component;
component FJK74E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    SD : in std_logic);
end component;
component FJK78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    J4 : in std_logic;
    J5 : in std_logic;
    J6 : in std_logic;
    J7 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    K4 : in std_logic;
    K5 : in std_logic;
    K6 : in std_logic;
    K7 : in std_logic;
    SD : in std_logic);
end component;
component FJK78E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    J4 : in std_logic;
    J5 : in std_logic;
    J6 : in std_logic;
    J7 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    K4 : in std_logic;
    K5 : in std_logic;
    K6 : in std_logic;
    K7 : in std_logic;
    SD : in std_logic);
end component;
component FT11
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FT21
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component IB11
  port (
    Z0 : out std_logic;
    XI0 : in std_logic);
end component;
component ID11
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    CLK : in std_logic);
end component;
component ID11E
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic);
end component;
component ID14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    CLK : in std_logic);
end component;
component ID14E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    CLK : in std_logic);
end component;
component ID21
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    CLK : in std_logic);
end component;
component ID24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    CLK : in std_logic);
end component;
component ID28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    CLK : in std_logic);
end component;
component ID31
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    XI0 : in std_logic);
end component;
component ID31E
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic);
end component;
component ID34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID34E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID41
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID41E
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID44E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID51
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID51E
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID54E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IL11
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    G : in std_logic);
end component;
component IL14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    G : in std_logic);
end component;
component IL18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    G : in std_logic);
end component;
component IL21
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    G : in std_logic);
end component;
component IL24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    G : in std_logic);
end component;
component IL28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    G : in std_logic);
end component;
component IL31
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    XI0 : in std_logic);
end component;
component IL34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IL41
  port (
    Q0 : out std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component IL44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IL51
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component IL54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IT14
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;

component IT18
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    O4 : out std_logic;
    O5 : out std_logic;
    O6 : out std_logic;
    O7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component IT21
  port (
    O0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component IT24
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component IT28
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    O4 : out std_logic;
    O5 : out std_logic;
    O6 : out std_logic;
    O7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component LD11
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component LD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component LD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic);
end component;
component LD21
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    CD : in std_logic);
end component;
component LD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    CD : in std_logic);
end component;
component LD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    CD : in std_logic);
end component;
component LD31
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    PD : in std_logic);
end component;
component LD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    PD : in std_logic);
end component;
component LD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    PD : in std_logic);
end component;
component LD41
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD51
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD61
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    TG : in std_logic);
end component;
component LD64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    TG : in std_logic);
end component;
component LD68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    TG : in std_logic);
end component;
component LD71
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD81
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    TG : in std_logic);
end component;
component LD84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    TG : in std_logic);
end component;
component LD88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    TG : in std_logic);
end component;
component LD91
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD98
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDA1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDA8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDI14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component LDI18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic);
end component;
component LDI24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component LDI28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic);
end component;
component LDI34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LDI38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LDI44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LDI48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LSR1
  port (
    Q0 : out std_logic;
    S0 : in std_logic;
    R0 : in std_logic);
end component;
component LSR2
  port (
    Q0 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    R0 : in std_logic;
    R1 : in std_logic);
end component;
component MAG2
  port (
    GT : out std_logic;
    EQ : out std_logic;
    LT : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    GTI : in std_logic;
    EQI : in std_logic;
    LTI : in std_logic);
end component;
component MAG4
  port (
    GT : out std_logic;
    EQ : out std_logic;
    LT : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    GTI : in std_logic;
    EQI : in std_logic;
    LTI : in std_logic);
end component;
component MAG8
  port (
    GT : out std_logic;
    EQ : out std_logic;
    LT : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    GTI : in std_logic;
    EQI : in std_logic;
    LTI : in std_logic);
end component;
component MULT24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component MULT44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component MUX16
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic);
end component;
component MUX16E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic);
end component;
component MUX2
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    S0 : in std_logic);
end component;
component MUX22
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    S0 : in std_logic);
end component;
component MUX22E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX24E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX2E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX4
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX42
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    S0 : in std_logic);
end component;
component MUX42E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX44A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX44AE
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX44E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX4E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX8
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic);
end component;
component MUX82
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    S0 : in std_logic);
end component;
component MUX82E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX8E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic);
end component;
component OB11
  port (
    XO0 : out std_logic;
    A0 : in std_logic);
end component;
component OB21
  port (
    XO0 : out std_logic;
    A0 : in std_logic);
end component;
component OB24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic);
end component;
component OB28
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic);
end component;
component OD11
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic);
end component;
component OD11E
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic);
end component;
component OD14
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic);
end component;
component OD14E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component OD21
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic);
end component;
component OD24
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic);
end component;
component OD31
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic);
end component;
component OD31E
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic);
end component;
component OD34
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic);
end component;
component OD34E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component OD41
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    SD : in std_logic);
end component;
component OD41E
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component OD44
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component OD44E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component OD51
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    SD : in std_logic);
end component;
component OD51E
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component OD54
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component OD54E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component ODT11
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component ODT11E
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT14
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component ODT14E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT21
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component ODT21E
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component ODT24E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT31
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT31E
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT34
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT34E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT41
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT41E
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT44
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT44E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OL11
  port (
    XQ0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component OL14
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component OL21
  port (
    XQ0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component OL24
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component OL31
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component OL34
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component OL41
  port (
    XQ0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OL44
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OL51
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OL54
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OLT11
  port (
    XO0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT14
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT21
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT31
  port (
    XO0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OLT34
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OLT41
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OLT44
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OT11
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT14
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT18
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component OT21
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT28
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component OT31
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT34
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT38
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component OT41
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT44
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT48
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component PG1
  port (
    PGO1 : out std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PG2
  port (
    PGO2 : out std_logic;
    GI2 : in std_logic;
    PI2 : in std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PG3
  port (
    PGO3 : out std_logic;
    GI3 : in std_logic;
    PI3 : in std_logic;
    GI2 : in std_logic;
    PI2 : in std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PG4
  port (
    PGO4 : out std_logic;
    GI4 : in std_logic;
    PI4 : in std_logic;
    GI3 : in std_logic;
    PI3 : in std_logic;
    GI2 : in std_logic;
    PI2 : in std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PREN10
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic);
end component;
component PREN10E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic;
    EN : in std_logic);
end component;
component PREN16
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic;
    S9 : in std_logic;
    S10 : in std_logic;
    S11 : in std_logic;
    S12 : in std_logic;
    S13 : in std_logic;
    S14 : in std_logic);
end component;
component PREN16E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic;
    S9 : in std_logic;
    S10 : in std_logic;
    S11 : in std_logic;
    S12 : in std_logic;
    S13 : in std_logic;
    S14 : in std_logic;
    EN : in std_logic);
end component;
component PREN8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic);
end component;
component PREN8E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    EN : in std_logic);
end component;
component SRR11
  port (
    Q0 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component SRR14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component SRR18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component SRR21
  port (
    Q0 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR31
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR41
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component SRR44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component SRR48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component SRR51
  port (
    Q0 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component SRR54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component SRR58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component SRRL1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CAIR : in std_logic;
    CAIL : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    RL : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component SRRL1S
  port (
    Q0 : out std_logic;
    CAIL : in std_logic;
    CAIR : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    PS : in std_logic;
    RL : in std_logic;
    SD : in std_logic);
end component;
component SRRL4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAIR : in std_logic;
    CAIL : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    RL : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component SRRL4S
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAIL : in std_logic;
    CAIR : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    PS : in std_logic;
    RL : in std_logic;
    SD : in std_logic);
end component;
component SRRL8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAIR : in std_logic;
    CAIL : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    RL : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component SRRL8S
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAIL : in std_logic;
    CAIR : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    PS : in std_logic;
    RL : in std_logic;
    SD : in std_logic);
end component;
component SUBF1
  port (
    Z0 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic;
    BI : in std_logic);
end component;
component SUBF16A
  port (
    BO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic;
    BI : in std_logic);
end component;
component SUBF2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    BI : in std_logic);
end component;
component SUBF4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    BI : in std_logic);
end component;
component SUBF8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    BI : in std_logic);
end component;
component SUBF8A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    BI : in std_logic);
end component;
component SUBH1
  port (
    Z0 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic);
end component;
component SUBH16A
  port (
    BO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic);
end component;
component SUBH2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic);
end component;
component SUBH3
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic);
end component;
component SUBH4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component SUBH8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component SUBH8A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component TCVRDC
  port (
    A : inout std_logic;
    B : inout std_logic;
    ENA : in std_logic;
    ENB : in std_logic);
end component;
component TCVRSC
  port (
    A : inout std_logic;
    B : inout std_logic;
    EN : in std_logic);
end component;
component LVPECLIN
   port(
      P_IN                       :	in    STD_ULOGIC;
      N_IN                       :	in    STD_ULOGIC;
      O                          :	out   STD_ULOGIC);
end component;
component LVPECLOUT
   port(
      I                          :	in    STD_ULOGIC;
      P_OUT                      :	out   STD_ULOGIC;
      N_OUT                      :	out   STD_ULOGIC);
end component;
component LVPECLTRI
   port(
      I                          :	in    STD_ULOGIC;
      OE                         :	in    STD_ULOGIC;
      P_OUT                      :	out   STD_ULOGIC;
      N_OUT                      :	out   STD_ULOGIC);
end component;


component SPLL
   generic (in_freq : string;
            CLK_OUT_TO_PIN: STRING := "OFF";
            WAKE_ON_LOCK: STRING := "OFF");
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC);
end component;
component STDPLL
   generic (in_freq  : string  := "100.0";
            mult     : string  := "1";
            div      : string  := "1";
            post     : string  := "1";
            secdiv   : string  := "1";
            lock_cyc : integer := 1;
            CLK_OUT_TO_PIN: STRING := "OFF";
            WAKE_ON_LOCK: STRING := "OFF";
            pll_dly  : string  := "0.0");
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC;
      PLL_LOCK                       :	out   STD_ULOGIC);
end component;
component STDPLLX
   generic (in_freq  : string  := "100.0";
            mult     : string  := "1";
            div      : string  := "1";
            post     : string  := "1";
            secdiv   : string  := "1";
            CLK_OUT_TO_PIN: STRING := "OFF";
            WAKE_ON_LOCK: STRING := "OFF";
            lock_cyc : integer := 1;
            pll_dly  : string  := "0.0");
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      PLL_FBK                        :	in    STD_ULOGIC;
      PLL_RST                        :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC;
      SEC_OUT                        :	out   STD_ULOGIC;
      PLL_LOCK                       :	out   STD_ULOGIC);
end component;
component LVDSIN
   port(
      P_IN                           :	in    STD_ULOGIC;
      N_IN                           :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;
component BLVDSIN
   port(
      P_IN                           :	in    STD_ULOGIC;
      N_IN                           :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;
component LVDSOUT
   port(
      I                              :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component BLVDSOUT
   port(
      I                              :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component LVDSTRI
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component BLVDSTRI
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component LVDSIO
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_IO                           :	inout   STD_ULOGIC;
      N_IO                           :	inout   STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;
component BLVDSIO
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_IO                           :	inout   STD_ULOGIC;
      N_IO                           :	inout   STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;

end VHD_PKG;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE STD.TEXTIO.ALL;

package components is
constant DefaultTimingChecksOn : Boolean := True;
constant DefaultXon : Boolean := True;
constant DefaultMsgOn : Boolean := True;

function Str2int( L : string) return integer;
function Str2real( L : string) return REAL;

component SPLL
   generic (in_freq : string;
            CLK_OUT_TO_PIN: STRING := "OFF";
            WAKE_ON_LOCK: STRING := "OFF");
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC);
end component;
component STDPLL
   generic (in_freq  : string  := "100.0";
            mult     : string  := "1";
            div      : string  := "1";
            post     : string  := "1";
            secdiv   : string  := "1";
            CLK_OUT_TO_PIN: STRING := "OFF";
            WAKE_ON_LOCK: STRING := "OFF";
            lock_cyc : integer := 1;
            pll_dly  : string  := "0.0");
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC;
      PLL_LOCK                       :	out   STD_ULOGIC);
end component;
component STDPLLX
   generic (in_freq  : string  := "100.0";
            mult     : string  := "1";
            div      : string  := "1";
            post     : string  := "1";
            secdiv   : string  := "1";
            CLK_OUT_TO_PIN: STRING := "OFF";
            WAKE_ON_LOCK: STRING := "OFF";
            lock_cyc : integer := 1;
            pll_dly  : string  := "1");
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      PLL_FBK                        :	in    STD_ULOGIC;
      PLL_RST                        :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC;
      SEC_OUT                        :	out   STD_ULOGIC;
      PLL_LOCK                       :	out   STD_ULOGIC);
end component;
component LVDSIN
   port(
      P_IN                           :	in    STD_ULOGIC;
      N_IN                           :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;
component BLVDSIN
   port(
      P_IN                           :	in    STD_ULOGIC;
      N_IN                           :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;
component LVDSOUT
   port(
      I                              :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component BLVDSOUT
   port(
      I                              :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component LVDSTRI
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component BLVDSTRI
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
end component;
component LVDSIO
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_IO                           :	inout   STD_ULOGIC;
      N_IO                           :	inout   STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;
component BLVDSIO
   port(
      I                              :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_IO                           :	inout   STD_ULOGIC;
      N_IO                           :	inout   STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
end component;

component LVPECLIN
   port(
      P_IN                       :	in    STD_ULOGIC;
      N_IN                       :	in    STD_ULOGIC;
      O                          :	out   STD_ULOGIC);
end component;
component LVPECLOUT
   port(
      I                          :	in    STD_ULOGIC;
      P_OUT                      :	out   STD_ULOGIC;
      N_OUT                      :	out   STD_ULOGIC);
end component;
component LVPECLTRI
   port(
      I                          :	in    STD_ULOGIC;
      OE                         :	in    STD_ULOGIC;
      P_OUT                      :	out   STD_ULOGIC;
      N_OUT                      :	out   STD_ULOGIC);
end component;

	component SHFE 
		port( REF : IN std_logic;
			  DATA : IN std_logic);
	end component;

	component PW 
		port( PULSE : IN std_logic);
	end component;

	component INV 
		port( A0 : IN std_logic;
			  ZN0 : OUT std_logic);
	end component;

	component BUF 
		port( A0 : IN std_logic;
			  Z0 : OUT std_logic);
	end component;

	component LXOR2
		port(A0 : IN std_logic;
			 A1 : IN std_logic;
			 Z0 : OUT std_logic);
	end component;

	component FD11
		port(D0 : IN std_logic;
			 CLK : IN std_logic;
			 Q0 : OUT std_logic);
	end component;

	component FD21
		port(D0 : IN std_logic;
			 CLK : IN std_logic;
			 CD : IN std_logic;
			 Q0 : OUT std_logic);
	end component;

	component XINV 
		port( A0 : IN std_logic;
			  ZN0 : OUT std_logic);
	end component;

	component XINPUT 
		port( XI0 : IN std_logic;
			  Z0 : OUT std_logic);
	end component;

	component XOUTPUT 
		port( A0 : IN std_logic;
			  XO0 : OUT std_logic);
	end component;

	component XBIDI1 
		port ( A0 : IN std_logic;
			   OE : IN std_logic;
			   Z0 : OUT std_logic;
			   XB0 : INOUT std_logic);
	 end component;

	component XTRI1 
		port( A0 : IN  std_logic;
			  OE : IN  std_logic;
			  XO0 : OUT  std_logic);
	end component;

	component XDFF1
		port( D0 : IN std_logic;
			  CLK : IN std_logic;
			  Q0 : OUT std_logic);
	end component;

	component XDL1
		port ( D0 : IN std_logic;
				G : IN std_logic;
			   Q0 : OUT std_logic);
	end component;

component XOR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component XOR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component OR16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND13 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND14 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND15 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND17 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 A16 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component AND18 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 A16 : IN std_logic;
		 A17 : IN std_logic;
		 Z0 : OUT std_logic);

end component;

component NAND2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NAND16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR5 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR6 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR10 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR11 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR12 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component NOR16 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR2 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR3 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR4 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR7 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR8 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component XNOR9 
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end component;

component FD11E
  port (D0, CLK, EN : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component FD21E
  port (D0, CLK, CD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component FDC1
  port (D0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component FDC1E
  port (D0, CLK, SD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component FDE1
  port (D0, CLK, CD, SD : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component FDE1E
  port (D0, CLK, CD, SD, EN : IN std_logic;
	               Q0 : OUT std_logic);
end component;

component FTI21
  port (T0, CLK, CD : IN std_logic;
                 Q0 : OUT std_logic);
end component;

component FTI21E
  port (T0, CLK, CD, EN : IN std_logic;
                     Q0 : OUT std_logic);
end component;

component FTI31
  port (T0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component FTI31E
  port (T0, CLK, SD, EN : IN std_logic;
		 Q0 : OUT std_logic);
end component;

component FTI41
  port (T0, CLK, SD, CD : IN std_logic;
		 Q0 : OUT std_logic);
end component;

component FTI41E
  port (T0, CLK, CD, SD, EN : IN std_logic;
		     Q0 : OUT std_logic);
end component;

component IT11
  port(A0, OE : IN std_logic;
	 O0 : OUT  std_logic);
end component;
       
component LDI11
  port (D0, G : IN std_logic;
           Q0 : OUT std_logic);
end component;

component LDI21
  port (D0, G, CD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component LDI31
  port (D0, G, SD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component LDI41
  port (D0, G, CD, SD : IN std_logic;
	         Q0 : OUT std_logic);
end component;

component XDFF1E
  port (D0, CLK, EN : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component XDFF2
  port (D0, CLK, CD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component XDFF2E
  port (D0, CLK, CD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component XDFF3
  port (D0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end component;

component XDFF3E
  port (D0, CLK, SD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component XDFF4
  port (D0, CLK, CD, SD : IN std_logic;
	           Q0 : OUT std_logic);
end component;

component XDFF4E
  port (D0, CLK, CD, SD, EN : IN std_logic;
	               Q0 : OUT std_logic);
end component;

component XDL2
  port (D0, G, CD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component XDL3
  port (D0, G, SD : IN std_logic;
	     Q0 : OUT std_logic);
end component;

component XDL4
  port (D0, G, CD, SD : IN std_logic;
	         Q0 : OUT std_logic);
end component;

component ADDF1
  port (
    Z0 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic;
    CI : in std_logic);
end component;
component ADDF16A
  port (
    CO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic;
    CI : in std_logic);
end component;
component ADDF2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    CI : in std_logic);
end component;
component ADDF4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    CI : in std_logic);
end component;
component ADDF8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    CI : in std_logic);
end component;
component ADDF8A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    CI : in std_logic);
end component;
component ADDH1
  port (
    Z0 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic);
end component;
component ADDH16A
  port (
    CO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic);
end component;
component ADDH2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic);
end component;
component ADDH3
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic);
end component;
component ADDH4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component ADDH8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    CO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component ADDH8A
  port (
    CO : out std_logic;
    Z7 : out std_logic;
    Z6 : out std_logic;
    Z5 : out std_logic;
    Z4 : out std_logic;
    Z3 : out std_logic;
    Z2 : out std_logic;
    Z1 : out std_logic;
    Z0 : out std_logic;
    B7 : in std_logic;
    B6 : in std_logic;
    B5 : in std_logic;
    B4 : in std_logic;
    B3 : in std_logic;
    B2 : in std_logic;
    B1 : in std_logic;
    B0 : in std_logic;
    A7 : in std_logic;
    A6 : in std_logic;
    A5 : in std_logic;
    A4 : in std_logic;
    A3 : in std_logic;
    A2 : in std_logic;
    A1 : in std_logic;
    A0 : in std_logic);
end component;
component BI11
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI14
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI18
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BI21
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI28
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BI31
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI34
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI38
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BI41
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component BI44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component BI48
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component BIID11
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID11E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIID14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID14E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIID18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID21
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID31
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID41
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID51
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID61
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID71
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID81
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID91
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID91E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIID94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic);
end component;
component BIID94E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIIDA1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDA1E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDA4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB1E
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIDB4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIIL11
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL21
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL31
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL41
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL51
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL61
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL71
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL81
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    XB4 : inout std_logic;
    XB5 : inout std_logic;
    XB6 : inout std_logic;
    XB7 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL91
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIIL94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIILA1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIILA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIILB1
  port (
    Q0 : out std_logic;
    XB0 : inout std_logic;
    A0 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIILB4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    CD : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIN27
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic);
end component;
component BIOD11
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component BIOD11E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD14
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component BIOD14E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD21
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component BIOD21E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component BIOD24E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component BIOD31
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD31E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD34
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD34E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD41
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD41E
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOD44E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL11
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL14
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL21
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component BIOL31
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL34
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL41
  port (
    Z0 : out std_logic;
    XB0 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component BIOL44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    XB0 : inout std_logic;
    XB1 : inout std_logic;
    XB2 : inout std_logic;
    XB3 : inout std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component CBD11
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD12
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBD21
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD22
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD31
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD32
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD41
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD42
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBD516
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD616
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CAO : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBD84
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBD88
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBD94
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBD98
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBDA16
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D10 : in std_logic;
    D11 : in std_logic;
    D12 : in std_logic;
    D13 : in std_logic;
    D14 : in std_logic;
    D15 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    D8 : in std_logic;
    D9 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDA4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDA8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDB4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBDB8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBU11
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU12
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component CBU21
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU22
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU31
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU32
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU41
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU42
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CBU516
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU616
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    CAO : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CBU716
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D10 : in std_logic;
    D11 : in std_logic;
    D12 : in std_logic;
    D13 : in std_logic;
    D14 : in std_logic;
    D15 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    D8 : in std_logic;
    D9 : in std_logic;
    EN : in std_logic;
    LD : in std_logic);
end component;
component CBU84
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBU88
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBU94
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBU98
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component CBUA16
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q10 : out std_logic;
    Q11 : out std_logic;
    Q12 : out std_logic;
    Q13 : out std_logic;
    Q14 : out std_logic;
    Q15 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    Q8 : out std_logic;
    Q9 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D10 : in std_logic;
    D11 : in std_logic;
    D12 : in std_logic;
    D13 : in std_logic;
    D14 : in std_logic;
    D15 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    D8 : in std_logic;
    D9 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUA4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUA8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUB4
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUB8
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUD1
  port (
    Q0 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD2
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD4S
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    DNUP : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CBUD8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CBUD8S
  port (
    CAO : out std_logic;
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    DNUP : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CDD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CDU44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDU48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CDUD4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CDUD4C
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CDUD8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CDUD8C
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAO : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CGD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CGD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CGD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CGU14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component CGU24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component CGU34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CGUD4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    DNUP : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component CGUD4S
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    DNUP : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component CMP2
  port (
    EQ : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic);
end component;
component CMP4
  port (
    EQ : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component CMP8
  port (
    EQ : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component DEC2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    S0 : in std_logic);
end component;
component DEC2E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DEC3
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DEC3E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DEC4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DEC4E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX22
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX22E
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DMUX24
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX24E
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX2E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DMUX4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX42
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX42E
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component DMUX44
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    W2 : out std_logic;
    W3 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    X2 : out std_logic;
    X3 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX44E
  port (
    W0 : out std_logic;
    W1 : out std_logic;
    W2 : out std_logic;
    W3 : out std_logic;
    X0 : out std_logic;
    X1 : out std_logic;
    X2 : out std_logic;
    X3 : out std_logic;
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX4E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component DMUX82
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Y4 : out std_logic;
    Y5 : out std_logic;
    Y6 : out std_logic;
    Y7 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    S0 : in std_logic);
end component;
component DMUX82E
  port (
    Y0 : out std_logic;
    Y1 : out std_logic;
    Y2 : out std_logic;
    Y3 : out std_logic;
    Y4 : out std_logic;
    Y5 : out std_logic;
    Y6 : out std_logic;
    Y7 : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component F3ADD
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    G012 : out std_logic;
    P012 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    CI : in std_logic);
end component;
component F3SUB
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    G012 : out std_logic;
    P012 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    BI : in std_logic);
end component;
component FD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic);
end component;
component FD14E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component FD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic);
end component;
component FD18E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic);
end component;
component FD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FD24E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component FD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FD28E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic);
end component;
component FD31
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic);
end component;
component FD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic);
end component;
component FD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic);
end component;
component FD41
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FD51
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component FD54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component FD58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component FD61
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FD64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FD68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FD71
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD81
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    TE : in std_logic);
end component;
component FD84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    TE : in std_logic);
end component;
component FD88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    TE : in std_logic);
end component;
component FD91
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FD98
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FDA1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic;
    TE : in std_logic);
end component;
component FDA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic;
    TE : in std_logic);
end component;
component FDA8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic;
    TE : in std_logic);
end component;
component FDB1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    SD : in std_logic);
end component;
component FDB4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CLK : in std_logic;
    SD : in std_logic);
end component;
component FDB8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CLK : in std_logic;
    SD : in std_logic);
end component;
component FDC4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component FDC4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FDC8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    SD : in std_logic);
end component;
component FDC8E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FDE4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component FDE4E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FDE8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    SD : in std_logic);
end component;
component FDE8E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component FJK11
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    CLK : in std_logic);
end component;
component FJK21
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FJK31
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    TE : in std_logic);
end component;
component FJK41
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    TI0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic;
    TE : in std_logic);
end component;
component FJK51
  port (
    Q0 : out std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CD : in std_logic);
end component;
component FJK61
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    SD : in std_logic);
end component;
component FJK64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    SD : in std_logic);
end component;
component FJK68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    J4 : in std_logic;
    J5 : in std_logic;
    J6 : in std_logic;
    J7 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    K4 : in std_logic;
    K5 : in std_logic;
    K6 : in std_logic;
    K7 : in std_logic;
    SD : in std_logic);
end component;
component FJK71
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    SD : in std_logic);
end component;
component FJK71E
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    J0 : in std_logic;
    K0 : in std_logic;
    SD : in std_logic);
end component;
component FJK74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    SD : in std_logic);
end component;
component FJK74E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    SD : in std_logic);
end component;
component FJK78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    J4 : in std_logic;
    J5 : in std_logic;
    J6 : in std_logic;
    J7 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    K4 : in std_logic;
    K5 : in std_logic;
    K6 : in std_logic;
    K7 : in std_logic;
    SD : in std_logic);
end component;
component FJK78E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    J0 : in std_logic;
    J1 : in std_logic;
    J2 : in std_logic;
    J3 : in std_logic;
    J4 : in std_logic;
    J5 : in std_logic;
    J6 : in std_logic;
    J7 : in std_logic;
    K0 : in std_logic;
    K1 : in std_logic;
    K2 : in std_logic;
    K3 : in std_logic;
    K4 : in std_logic;
    K5 : in std_logic;
    K6 : in std_logic;
    K7 : in std_logic;
    SD : in std_logic);
end component;
component FT11
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component FT21
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    CS : in std_logic);
end component;
component IB11
  port (
    Z0 : out std_logic;
    XI0 : in std_logic);
end component;
component ID11
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    CLK : in std_logic);
end component;
component ID11E
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic);
end component;
component ID14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    CLK : in std_logic);
end component;
component ID14E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    CLK : in std_logic);
end component;
component ID21
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    CLK : in std_logic);
end component;
component ID24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    CLK : in std_logic);
end component;
component ID28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    CLK : in std_logic);
end component;
component ID31
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    XI0 : in std_logic);
end component;
component ID31E
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic);
end component;
component ID34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID34E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID41
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID41E
  port (
    Q0 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID44E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID51
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID51E
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component ID54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component ID54E
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IL11
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    G : in std_logic);
end component;
component IL14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    G : in std_logic);
end component;
component IL18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    G : in std_logic);
end component;
component IL21
  port (
    Q0 : out std_logic;
    XI0 : in std_logic;
    G : in std_logic);
end component;
component IL24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    G : in std_logic);
end component;
component IL28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic;
    XI4 : in std_logic;
    XI5 : in std_logic;
    XI6 : in std_logic;
    XI7 : in std_logic;
    G : in std_logic);
end component;
component IL31
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    XI0 : in std_logic);
end component;
component IL34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IL41
  port (
    Q0 : out std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component IL44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IL51
  port (
    Q0 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic);
end component;
component IL54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    G : in std_logic;
    SD : in std_logic;
    XI0 : in std_logic;
    XI1 : in std_logic;
    XI2 : in std_logic;
    XI3 : in std_logic);
end component;
component IT14
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;

component IT18
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    O4 : out std_logic;
    O5 : out std_logic;
    O6 : out std_logic;
    O7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component IT21
  port (
    O0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component IT24
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component IT28
  port (
    O0 : out std_logic;
    O1 : out std_logic;
    O2 : out std_logic;
    O3 : out std_logic;
    O4 : out std_logic;
    O5 : out std_logic;
    O6 : out std_logic;
    O7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component LD11
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component LD14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component LD18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic);
end component;
component LD21
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    CD : in std_logic);
end component;
component LD24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    CD : in std_logic);
end component;
component LD28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    CD : in std_logic);
end component;
component LD31
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    PD : in std_logic);
end component;
component LD34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    PD : in std_logic);
end component;
component LD38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    PD : in std_logic);
end component;
component LD41
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD51
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic);
end component;
component LD61
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    TG : in std_logic);
end component;
component LD64
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    TG : in std_logic);
end component;
component LD68
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    TG : in std_logic);
end component;
component LD71
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD74
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD78
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD81
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    TG : in std_logic);
end component;
component LD84
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    TG : in std_logic);
end component;
component LD88
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    TG : in std_logic);
end component;
component LD91
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD94
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LD98
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDA1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    TI0 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDA4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDA8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    TI0 : in std_logic;
    TI1 : in std_logic;
    TI2 : in std_logic;
    TI3 : in std_logic;
    TI4 : in std_logic;
    TI5 : in std_logic;
    TI6 : in std_logic;
    TI7 : in std_logic;
    G : in std_logic;
    PD : in std_logic;
    CD : in std_logic;
    TG : in std_logic);
end component;
component LDI14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component LDI18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic);
end component;
component LDI24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component LDI28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic);
end component;
component LDI34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LDI38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LDI44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LDI48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component LSR1
  port (
    Q0 : out std_logic;
    S0 : in std_logic;
    R0 : in std_logic);
end component;
component LSR2
  port (
    Q0 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    R0 : in std_logic;
    R1 : in std_logic);
end component;
component MAG2
  port (
    GT : out std_logic;
    EQ : out std_logic;
    LT : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    GTI : in std_logic;
    EQI : in std_logic;
    LTI : in std_logic);
end component;
component MAG4
  port (
    GT : out std_logic;
    EQ : out std_logic;
    LT : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    GTI : in std_logic;
    EQI : in std_logic;
    LTI : in std_logic);
end component;
component MAG8
  port (
    GT : out std_logic;
    EQ : out std_logic;
    LT : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    GTI : in std_logic;
    EQI : in std_logic;
    LTI : in std_logic);
end component;
component MULT24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component MULT44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component MUX16
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic);
end component;
component MUX16E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic);
end component;
component MUX2
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    S0 : in std_logic);
end component;
component MUX22
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    S0 : in std_logic);
end component;
component MUX22E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX24
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX24E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX2E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX4
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX42
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    S0 : in std_logic);
end component;
component MUX42E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX44
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX44A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX44AE
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX44E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    C0 : in std_logic;
    C1 : in std_logic;
    C2 : in std_logic;
    C3 : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX4E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic);
end component;
component MUX8
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic);
end component;
component MUX82
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    S0 : in std_logic);
end component;
component MUX82E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic);
end component;
component MUX8E
  port (
    Z0 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    EN : in std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic);
end component;
component OB11
  port (
    XO0 : out std_logic;
    A0 : in std_logic);
end component;
component OB21
  port (
    XO0 : out std_logic;
    A0 : in std_logic);
end component;
component OB24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic);
end component;
component OB28
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic);
end component;
component OD11
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic);
end component;
component OD11E
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic);
end component;
component OD14
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic);
end component;
component OD14E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component OD21
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic);
end component;
component OD24
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic);
end component;
component OD31
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic);
end component;
component OD31E
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic);
end component;
component OD34
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic);
end component;
component OD34E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic);
end component;
component OD41
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    SD : in std_logic);
end component;
component OD41E
  port (
    XQ0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component OD44
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component OD44E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component OD51
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    SD : in std_logic);
end component;
component OD51E
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component OD54
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    SD : in std_logic);
end component;
component OD54E
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    SD : in std_logic);
end component;
component ODT11
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component ODT11E
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT14
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component ODT14E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT21
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic);
end component;
component ODT21E
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic);
end component;
component ODT24E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic);
end component;
component ODT31
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT31E
  port (
    XO0 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT34
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT34E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT41
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT41E
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT44
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component ODT44E
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OL11
  port (
    XQ0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component OL14
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component OL21
  port (
    XQ0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component OL24
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component OL31
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic);
end component;
component OL34
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic);
end component;
component OL41
  port (
    XQ0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OL44
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OL51
  port (
    XQ0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OL54
  port (
    XQ0 : out std_logic;
    XQ1 : out std_logic;
    XQ2 : out std_logic;
    XQ3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    SD : in std_logic);
end component;
component OLT11
  port (
    XO0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT14
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT21
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic);
end component;
component OLT31
  port (
    XO0 : out std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OLT34
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OLT41
  port (
    XO0 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OLT44
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    CD : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    G : in std_logic;
    OE : in std_logic;
    SD : in std_logic);
end component;
component OT11
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT14
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT18
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component OT21
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT24
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT28
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component OT31
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT34
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT38
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component OT41
  port (
    XO0 : out std_logic;
    A0 : in std_logic;
    OE : in std_logic);
end component;
component OT44
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    OE : in std_logic);
end component;
component OT48
  port (
    XO0 : out std_logic;
    XO1 : out std_logic;
    XO2 : out std_logic;
    XO3 : out std_logic;
    XO4 : out std_logic;
    XO5 : out std_logic;
    XO6 : out std_logic;
    XO7 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    OE : in std_logic);
end component;
component PG1
  port (
    PGO1 : out std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PG2
  port (
    PGO2 : out std_logic;
    GI2 : in std_logic;
    PI2 : in std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PG3
  port (
    PGO3 : out std_logic;
    GI3 : in std_logic;
    PI3 : in std_logic;
    GI2 : in std_logic;
    PI2 : in std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PG4
  port (
    PGO4 : out std_logic;
    GI4 : in std_logic;
    PI4 : in std_logic;
    GI3 : in std_logic;
    PI3 : in std_logic;
    GI2 : in std_logic;
    PI2 : in std_logic;
    GI1 : in std_logic;
    PI1 : in std_logic;
    PGI1 : in std_logic);
end component;
component PREN10
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic);
end component;
component PREN10E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic;
    EN : in std_logic);
end component;
component PREN16
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic;
    S9 : in std_logic;
    S10 : in std_logic;
    S11 : in std_logic;
    S12 : in std_logic;
    S13 : in std_logic;
    S14 : in std_logic);
end component;
component PREN16E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    S7 : in std_logic;
    S8 : in std_logic;
    S9 : in std_logic;
    S10 : in std_logic;
    S11 : in std_logic;
    S12 : in std_logic;
    S13 : in std_logic;
    S14 : in std_logic;
    EN : in std_logic);
end component;
component PREN8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic);
end component;
component PREN8E
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    S0 : in std_logic;
    S1 : in std_logic;
    S2 : in std_logic;
    S3 : in std_logic;
    S4 : in std_logic;
    S5 : in std_logic;
    S6 : in std_logic;
    EN : in std_logic);
end component;
component SRR11
  port (
    Q0 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component SRR14
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component SRR18
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    CD : in std_logic);
end component;
component SRR21
  port (
    Q0 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR24
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR28
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR31
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR34
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR38
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CD : in std_logic);
end component;
component SRR41
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component SRR44
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component SRR48
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAI : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    CS : in std_logic);
end component;
component SRR51
  port (
    Q0 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component SRR54
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component SRR58
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAI : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    SD : in std_logic);
end component;
component SRRL1
  port (
    Q0 : out std_logic;
    D0 : in std_logic;
    CAIR : in std_logic;
    CAIL : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    RL : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component SRRL1S
  port (
    Q0 : out std_logic;
    CAIL : in std_logic;
    CAIR : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    PS : in std_logic;
    RL : in std_logic;
    SD : in std_logic);
end component;
component SRRL4
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    CAIR : in std_logic;
    CAIL : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    RL : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component SRRL4S
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    CAIL : in std_logic;
    CAIR : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    PS : in std_logic;
    RL : in std_logic;
    SD : in std_logic);
end component;
component SRRL8
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    CAIR : in std_logic;
    CAIL : in std_logic;
    CLK : in std_logic;
    PS : in std_logic;
    LD : in std_logic;
    EN : in std_logic;
    RL : in std_logic;
    CD : in std_logic;
    CS : in std_logic);
end component;
component SRRL8S
  port (
    Q0 : out std_logic;
    Q1 : out std_logic;
    Q2 : out std_logic;
    Q3 : out std_logic;
    Q4 : out std_logic;
    Q5 : out std_logic;
    Q6 : out std_logic;
    Q7 : out std_logic;
    CAIL : in std_logic;
    CAIR : in std_logic;
    CD : in std_logic;
    CLK : in std_logic;
    CS : in std_logic;
    D0 : in std_logic;
    D1 : in std_logic;
    D2 : in std_logic;
    D3 : in std_logic;
    D4 : in std_logic;
    D5 : in std_logic;
    D6 : in std_logic;
    D7 : in std_logic;
    EN : in std_logic;
    LD : in std_logic;
    PS : in std_logic;
    RL : in std_logic;
    SD : in std_logic);
end component;
component SUBF1
  port (
    Z0 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic;
    BI : in std_logic);
end component;
component SUBF16A
  port (
    BO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic;
    BI : in std_logic);
end component;
component SUBF2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    BI : in std_logic);
end component;
component SUBF4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    BI : in std_logic);
end component;
component SUBF8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    BI : in std_logic);
end component;
component SUBF8A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    BI : in std_logic);
end component;
component SUBH1
  port (
    Z0 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    B0 : in std_logic);
end component;
component SUBH16A
  port (
    BO : out std_logic;
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z10 : out std_logic;
    Z11 : out std_logic;
    Z12 : out std_logic;
    Z13 : out std_logic;
    Z14 : out std_logic;
    Z15 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    Z8 : out std_logic;
    Z9 : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A10 : in std_logic;
    A11 : in std_logic;
    A12 : in std_logic;
    A13 : in std_logic;
    A14 : in std_logic;
    A15 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    A8 : in std_logic;
    A9 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B10 : in std_logic;
    B11 : in std_logic;
    B12 : in std_logic;
    B13 : in std_logic;
    B14 : in std_logic;
    B15 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic;
    B8 : in std_logic;
    B9 : in std_logic);
end component;
component SUBH2
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic);
end component;
component SUBH3
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic);
end component;
component SUBH4
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic);
end component;
component SUBH8
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component SUBH8A
  port (
    Z0 : out std_logic;
    Z1 : out std_logic;
    Z2 : out std_logic;
    Z3 : out std_logic;
    Z4 : out std_logic;
    Z5 : out std_logic;
    Z6 : out std_logic;
    Z7 : out std_logic;
    BO : out std_logic;
    A0 : in std_logic;
    A1 : in std_logic;
    A2 : in std_logic;
    A3 : in std_logic;
    A4 : in std_logic;
    A5 : in std_logic;
    A6 : in std_logic;
    A7 : in std_logic;
    B0 : in std_logic;
    B1 : in std_logic;
    B2 : in std_logic;
    B3 : in std_logic;
    B4 : in std_logic;
    B5 : in std_logic;
    B6 : in std_logic;
    B7 : in std_logic);
end component;
component TCVRDC
  port (
    A : inout std_logic;
    B : inout std_logic;
    ENA : in std_logic;
    ENB : in std_logic);
end component;
component TCVRSC
  port (
    A : inout std_logic;
    B : inout std_logic;
    EN : in std_logic);
end component;
end components;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.std_logic_arith.all;

package body components is 
 
 
 function str2int( L : string) return integer is
	variable ok:         boolean;
	variable pos:        integer:=1;
	variable sign: integer := 1;
	variable rval: integer := 0;
	variable value: integer := 0;
    begin
	ok := FALSE;
	if pos < L'right and (L(pos) = '-' or L(pos) = '+') then
	    if L(pos) = '-' then
		sign := -1;
	    end if;
	    pos := pos + 1;
	end if;

	-- Once the optional leading sign is removed, an integer can
	--   contain only the digits '0' through '9' and the '_'
	--   (underscore) character.  VHDL disallows two successive
	--   underscores, and leading or trailing underscores.

	if pos <= L'right and L(pos) >= '0' and L(pos) <= '9' then
	    while pos <= L'right loop
		if L(pos) >= '0' and L(pos) <= '9' then
		    rval := rval * 10
		            + character'pos(L(pos)) - character'pos('0');
		    ok := TRUE;
		elsif L(pos) = '_' then
		    if pos = L'right
		    or L(pos + 1) < '0'
		    or L(pos + 1) > '9' then
			ok := FALSE;
			exit;
		    end if;
		else
		    exit;
		end if;
		pos := pos + 1;
	    end loop;
	end if;

	value := sign * rval;
        RETURN(value);
    end str2int;

    function str2real( L: string) return real is
	variable pos:        integer;
	variable value:      real;
	variable value1:      real;
	variable ok:         boolean;
	variable sign:       real := 1.0;
	variable rval:       real := 0.0;
        variable powerten:   real := 0.1;

        begin

	pos := L'left;
	if (pos <= L'right) and (L(pos) = '-') then
	    sign := -1.0;
	    pos := pos + 1;
	end if;

            ok := FALSE;
            rval := 0.0;
            if pos <= L'right and L(pos) >= '0' and L(pos) <= '9' then
                while pos <= L'right and L(pos) /= '.' and L(pos) /= ' ' and L(pos) /= HT  loop
                    if L(pos) >= '0' and L(pos) <= '9' then
                        rval := rval*10.0 + real(character'pos(L(pos)) - character'pos('0'));
                        pos := pos+1;
                        ok := true;
                    else
                        ok := false;
                        exit;
                    end if;
                end loop;
            end if;

	    if ok and pos <= L'right and L(pos) = '.' then
	    pos := pos + 1;
            end if;

            if pos <= L'right then
               while pos <= L'right and ((L(pos) >= '0' and L(pos) <= '9') or L(pos) = '_') loop
                       rval := rval + (real(character'pos(L(pos))-character'pos('0'))*powerten);
                       powerten := powerten*0.1;
                      pos := pos+1;
                     ok := true;
            end loop;
        end if;

        if ok then
            value := rval * sign;
        end if;

        if (L'right <= 2) then
           value1 := 0.25 * value;
        else
           value1 := value;
        end if;

        return (value1);
      end str2real;
 
end components;


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library lat_vhd;
use lat_vhd.components.all;


-- entity declaration --
entity SPLL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      IN_FREQ: STRING := "100.0";
      CLK_OUT_TO_PIN: STRING := "OFF";
      WAKE_ON_LOCK: STRING := "OFF";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_IN_CLK_OUT             :	VitalDelayType01 := (0.00 ns, 0.00 ns);
      tipd_CLK_IN                    :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      CLK_IN                         :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of SPLL : entity is FALSE;
end SPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of SPLL is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL CLK_IN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (CLK_IN_ipd, CLK_IN, tipd_CLK_IN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (CLK_IN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(CLK_IN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CLK_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "CLK_OUT",
       OutTemp => O_zd,
       Paths => (0 => (CLK_IN_ipd'last_event, tpd_CLK_IN_CLK_OUT, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell STDPLL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library lattice;
use lattice.components.all;

-- entity declaration --
entity STDPLL is
   generic(
      IN_FREQ  : string  := "100.0";
      CLK_OUT_TO_PIN: STRING := "OFF";
      WAKE_ON_LOCK: STRING := "OFF";
      MULT     : string  := "1";
      DIV      : string  := "1";
      POST     : string  := "1";
      SECDIV   : string  := "2";
      lock_cyc : integer := 2;
      PLL_DLY  : string  := "0.0";
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_CLK_IN_CLK_OUT             :	VitalDelayType01 := (0.00 ns, 0.00 ns);
      tpd_CLK_IN_PLL_LOCK             :	VitalDelayType01 := (0.00 ns, 0.00 ns);
      tipd_CLK_IN             :	VitalDelayType01 := (0.000 ns, 0.000 ns));
   port(
      CLK_IN                         :	in    STD_ULOGIC;
      CLK_OUT                        :	out   STD_ULOGIC;
      PLL_LOCK                       :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of STDPLL : entity is FALSE;
end STDPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library lattice;
use lattice.components.all;
architecture VITAL of STDPLL is
   attribute VITAL_LEVEL1 of VITAL : architecture is FALSE;

   SIGNAL CLK_IN_ipd	 : STD_ULOGIC := 'X';

  CONSTANT input_frequency : REAL := str2real(in_freq);

  SIGNAL clklock_half_period : TIME :=100 ns;
  SIGNAL clklock_half_period1 : TIME :=100 ns;
  SIGNAL clklock_half_period0 : TIME :=100 ns;
  SIGNAL clklock_half_period_minus_dly1 : TIME :=100 ns;
  SIGNAL clklock_half_period_minus_dly0 : TIME :=100 ns;
  SIGNAL start_inclk : STD_LOGIC ;
  SIGNAL clklock_rising_edge_count : INTEGER := 0 ;
  SIGNAL clklock_falling_edge_count : INTEGER := 0 ;
  SIGNAL clklock_last_rising_edge : TIME ;
  SIGNAL clklock_last_falling_edge : TIME ;

  SIGNAL clock_count : INTEGER := -1 ;
  SIGNAL clklock_lock : BOOLEAN := TRUE;
  SIGNAL CLK_OUT_sig_d  : std_logic := '0';
  SIGNAL CLK_OUT_sig_d_not  : std_logic := '0';
  SIGNAL CLK_OUT_start  : std_logic := '0';
  SIGNAL CLK_OUT_sig_3d  : std_logic := '0';
  SIGNAL CLK_OUT_sig_d_start  : std_logic := '0';
  SIGNAL CLK_OUT_sig1 : std_logic := '0';
  SIGNAL CLK_OUT_plus_delay : std_logic := '0';
  SIGNAL PLL_LOCK_plus : std_logic := '0';
  SIGNAL PLL_LOCK_minus : std_logic := '0';
  CONSTANT clockboost: integer := str2int(mult) / str2int(div);
  CONSTANT tpd: time := 1.0 ns * str2real(pll_dly);

BEGIN

   WireDelay : block
   begin
   VitalWireDelay (CLK_IN_ipd, CLK_IN, tipd_CLK_IN);
   end block;

edge_count: PROCESS
     VARIABLE input_cycle : REAL;
     VARIABLE real_cycle : REAL;
BEGIN
     clklock_half_period <= (clklock_half_period0 + clklock_half_period1)/2;

  WAIT UNTIL (CLK_IN_ipd'EVENT AND CLK_IN_ipd='1');	   
     clklock_rising_edge_count <= clklock_rising_edge_count +1;
     IF clklock_rising_edge_count = 0 THEN
        clklock_last_rising_edge <= NOW;	
	start_inclk <= CLK_IN_ipd;
     ELSE
     IF clklock_rising_edge_count = 1 THEN
       clklock_half_period0 <= (NOW - clklock_last_falling_edge)* real(str2int(div))/real(str2int(mult));
	input_cycle := 1000.0 / input_frequency;
	real_cycle := REAL( (NOW - clklock_last_rising_edge) / 1 ns);
	IF ( real_cycle < 0.9 * input_cycle OR
	     real_cycle > 1.1 * input_cycle ) THEN
  	      	ASSERT TRUE 
  		REPORT " Input_Frequency Violation "
  		SEVERITY WARNING;
  		clklock_lock <= FALSE;
        END IF;
       clklock_half_period_minus_dly0 <= (NOW - clklock_last_falling_edge) + tpd;
     END IF;
     END IF;
 
  WAIT UNTIL (CLK_IN_ipd'EVENT AND CLK_IN_ipd='0');
     clklock_falling_edge_count <= clklock_falling_edge_count +1;	  	
     IF clklock_falling_edge_count = 0 THEN	
	clklock_last_falling_edge <= NOW;
	clklock_half_period1 <= (NOW - clklock_last_rising_edge)* real(str2int(div))/real(str2int(mult)); 
     ELSIF clklock_falling_edge_count = 1 THEN
        clklock_half_period_minus_dly1 <= (NOW - clklock_last_rising_edge) + tpd;
     END IF;
END PROCESS edge_count;

toggle: PROCESS
BEGIN

     WAIT ON clklock_rising_edge_count;
     IF clklock_rising_edge_count > lock_cyc + 1 THEN
        if(clockboost >1) then
	   FOR i IN 1 TO (2*clockboost) LOOP 	         
		clock_count <= clock_count + 1;
		WAIT FOR clklock_half_period;
	END LOOP;
      else  
		clock_count <= clock_count + 1;
		WAIT FOR (clklock_half_period);
      end if;
     ELSE
	clock_count <= 0;
     END IF;
END PROCESS toggle;


gen_pll_lock_plus:process
begin
     wait until (clock_count=1);
          PLL_LOCK_plus <= '1';
end process;

gen_pll_lock_minus:process
begin
     wait until (clock_count=3);
          PLL_LOCK_minus <= '1';
end process;

process
begin 
    wait until clock_count = 1;
    CLK_OUT_sig_d_start <='1';
end process;

process
begin
   wait until CLK_OUT_sig_d_start = '1'; LOOP
     wait for clklock_half_period1;
   CLK_OUT_sig_d_not <= not CLK_OUT_sig_d_not;
     wait for clklock_half_period0;
   CLK_OUT_sig_d_not <= not CLK_OUT_sig_d_not ;
   END LOOP;
end process;

process(clklock_falling_edge_count)
begin
   if (clklock_falling_edge_count >= lock_cyc + 1) then
       CLK_OUT_start <= '1' after clklock_half_period_minus_dly0;
   end if;
end process;

process
begin
   wait until  CLK_OUT_start = '1'; LOOP
      CLK_OUT_sig_3d <= not CLK_OUT_sig_3d;
     wait for clklock_half_period1;
      CLK_OUT_sig_3d <= not CLK_OUT_sig_3d ;
     wait for clklock_half_period0;
     END LOOP;
end process;


    CLK_OUT_sig_d <= CLK_OUT_sig_d_start and not CLK_OUT_sig_d_not; 

    CLK_OUT_plus_delay <= CLK_OUT_sig_d after tpd when tpd >= 0 ns else
                          CLK_OUT_sig_3d; 

    CLK_OUT <= CLK_OUT_plus_delay;

    PLL_LOCK <= PLL_LOCK_plus when tpd >= 0 ns else
                PLL_LOCK_minus;
               

end VITAL;

configuration CFG_STDPLL_VITAL of STDPLL is 
        for VITAL
        end for; 
end CFG_STDPLL_VITAL;


----- VITAL model for cell STDPLLX -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;
library lattice;
use lattice.components.all;

-- entity declaration --
entity STDPLLX is
   generic(
      IN_FREQ  : string  := "100.0";
      CLK_OUT_TO_PIN: STRING := "OFF";
      WAKE_ON_LOCK: STRING := "OFF";
      MULT     : string  := "1";
      DIV      : string  := "1";
      POST     : string  := "1";
      LOCK_CYC : integer := 2;
      SECDIV   : string   := "2";
      PLL_DLY  : string  := "0.0";
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_PLL_RST_PLL_LOCK :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_CLK_IN_CLK_OUT             :	VitalDelayType01 := (0.00 ns, 0.00 ns);
      tpd_CLK_IN_PLL_LOCK             :	VitalDelayType01 := (0.00 ns, 0.00 ns);
      tpd_CLK_IN_SEC_OUT             :	VitalDelayType01 := (0.00 ns, 0.00 ns);
      tipd_CLK_IN             :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PLL_FBK   :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PLL_RST   :	VitalDelayType01 := (0.000 ns, 0.000 ns));
   port(
      CLK_IN            : in    STD_ULOGIC;
      PLL_FBK           : in    STD_ULOGIC;
      PLL_RST           : in    STD_ULOGIC;
      CLK_OUT           : out   STD_ULOGIC;
      SEC_OUT           : out   STD_ULOGIC;
      PLL_LOCK          : out   STD_ULOGIC);
attribute VITAL_LEVEL0 of STDPLLX : entity is FALSE;
end STDPLLX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library lattice;
use lattice.components.all;


architecture VITAL of STDPLLX is
  attribute VITAL_LEVEL1 of VITAL : architecture is FALSE;

  SIGNAL CLK_IN_ipd	 : STD_ULOGIC := 'X';
  SIGNAL PLL_RST_ipd	 : STD_ULOGIC := 'X';

  CONSTANT input_frequency : REAL := str2real(in_freq);

  SIGNAL clklock_half_period : TIME :=100 ns;
  SIGNAL clklock_half_period1 : TIME :=100 ns;
  SIGNAL clklock_half_period0 : TIME :=100 ns;
  SIGNAL clklock_half_period_minus_dly1 : TIME :=100 ns;
  SIGNAL clklock_half_period_minus_dly0 : TIME :=100 ns;
  SIGNAL secd_delay_minus1 : TIME :=100 ns;
  SIGNAL secd_delay_minus0 : TIME :=100 ns;
  SIGNAL start_inclk : STD_LOGIC ;
  SIGNAL clklock_rising_edge_count : INTEGER := 0 ;
  SIGNAL clklock_falling_edge_count : INTEGER := 0 ;
  SIGNAL clklock_last_rising_edge : TIME ;
  SIGNAL clklock_last_falling_edge : TIME ;

  SIGNAL clock_count : INTEGER := -1 ;
  SIGNAL clklock_lock : BOOLEAN := TRUE;
  SIGNAL CLK_OUT_sig_d  : std_logic := '0';
  SIGNAL CLK_OUT_sig_d_not  : std_logic := '0';

  SIGNAL CLK_OUT_sig_3d  : std_logic := '0';
  SIGNAL CLK_OUT_sig_d_start  : std_logic := '0';
  SIGNAL CLK_OUT_start  : std_logic := '0';
  SIGNAL CLK_OUT_plus_delay : std_logic := '0';
  SIGNAL SEC_OUT_sig_d  : std_logic := '0';
  SIGNAL SEC_OUT_sig_d_not  : std_logic := '0';

  SIGNAL SEC_OUT_sig_3d  : std_logic := '0';
  SIGNAL SEC_OUT_sig_d_start  : std_logic := '0';
  SIGNAL SEC_OUT_start  : std_logic := '0';
  SIGNAL SEC_OUT_plus_delay : std_logic := '0';
  SIGNAL CLK_OUT_sig1 : std_logic := '0';
  SIGNAL PLL_LOCK_plus : std_logic := '0';
  SIGNAL PLL_LOCK_minus : std_logic := '0';

  CONSTANT secdiv_p: integer := str2int(secdiv);
  CONSTANT clockboost: integer := str2int(mult) / str2int(div);
  CONSTANT tpd: time := 1.0 ns * str2real(pll_dly);

BEGIN
   WireDelay : block
   begin
   VitalWireDelay (CLK_IN_ipd, CLK_IN, tipd_CLK_IN);
   VitalWireDelay (PLL_RST_ipd, PLL_RST, tipd_PLL_RST);
   end block;

edge_count: PROCESS
     VARIABLE input_cycle : REAL;
     VARIABLE real_cycle : REAL;
BEGIN
      clklock_half_period <= (clklock_half_period0 + clklock_half_period1)/2;

  WAIT UNTIL (CLK_IN_ipd'EVENT AND CLK_IN_ipd='1');	   
     clklock_rising_edge_count <= clklock_rising_edge_count +1;
     IF clklock_rising_edge_count = 0 THEN
        clklock_last_rising_edge <= NOW;	
	start_inclk <= CLK_IN_ipd;
     ELSE
     IF clklock_rising_edge_count = 1 THEN
       clklock_half_period0 <= (NOW - clklock_last_falling_edge)* real(str2int(div))/real(str2int(mult));
	input_cycle := 1000.0 / input_frequency;
	real_cycle := REAL( (NOW - clklock_last_rising_edge) / 1 ns);
	IF ( real_cycle < 0.9 * input_cycle OR
	     real_cycle > 1.1 * input_cycle ) THEN
  	      	ASSERT TRUE 
  		REPORT " Input_Frequency Violation "
  		SEVERITY WARNING;
  		clklock_lock <= FALSE;
        END IF;
       clklock_half_period_minus_dly0 <= (NOW - clklock_last_falling_edge) + tpd;
        secd_delay_minus0 <= clklock_half_period0 * secdiv_p + tpd;
     END IF;
     END IF;
 
  WAIT UNTIL (CLK_IN_ipd'EVENT AND CLK_IN_ipd='0');
     clklock_falling_edge_count <= clklock_falling_edge_count +1;	  	
     IF clklock_falling_edge_count = 0 THEN	
	clklock_last_falling_edge <= NOW;
	clklock_half_period1 <= (NOW - clklock_last_rising_edge)* real(str2int(div))/real(str2int(mult)); 
     ELSIF clklock_falling_edge_count = 1 THEN
        clklock_half_period_minus_dly1 <= (NOW - clklock_last_rising_edge) + tpd;
        secd_delay_minus1 <= clklock_half_period1 * secdiv_p + tpd;
     END IF;
END PROCESS edge_count;

toggle: PROCESS
BEGIN

     WAIT ON clklock_rising_edge_count;
     IF clklock_rising_edge_count > lock_cyc + 1 and PLL_RST_ipd ='0' THEN
        if(clockboost >1) then
	   FOR i IN 1 TO (2*clockboost) LOOP 	       
		clock_count <= clock_count + 1;
		WAIT FOR clklock_half_period;
	   END LOOP;
        else  
		clock_count <= clock_count + 1;
		WAIT FOR (clklock_half_period);
        end if;
     ELSE
	clock_count <= 0;
     END IF;
END PROCESS toggle;


gen_pll_lock_plus:process
begin
     wait until (clock_count=1);
          PLL_LOCK_plus <= '1';
end process;

gen_pll_lock_minus:process
begin
     wait until (clock_count=3);
          PLL_LOCK_minus <= '1';
end process;

process
begin 
    wait until clock_count = 1;
    CLK_OUT_sig_d_start <='1';
    SEC_OUT_sig_d_start <='1';
end process;

process
begin
   wait until CLK_OUT_sig_d_start = '1'; LOOP
     wait for clklock_half_period1;
   CLK_OUT_sig_d_not <= not CLK_OUT_sig_d_not;
     wait for clklock_half_period0;
   CLK_OUT_sig_d_not <= not CLK_OUT_sig_d_not ;
   END LOOP;
end process;

process(clklock_falling_edge_count)
begin
   if (clklock_falling_edge_count >= lock_cyc + 1 and PLL_RST_ipd = '0') then
       CLK_OUT_start <= '1' after clklock_half_period_minus_dly0;
   end if;
end process;

process
begin
   wait until  CLK_OUT_start = '1'; LOOP
      CLK_OUT_sig_3d <= not CLK_OUT_sig_3d;
     wait for clklock_half_period1;
      CLK_OUT_sig_3d <= not CLK_OUT_sig_3d ;
     wait for clklock_half_period0;
     END LOOP;
end process;

process
begin
   wait until SEC_OUT_sig_d_start = '1'; LOOP
     wait for clklock_half_period1 * secdiv_p;
   SEC_OUT_sig_d_not <= not SEC_OUT_sig_d_not;
     wait for clklock_half_period0 * secdiv_p;
   SEC_OUT_sig_d_not <= not SEC_OUT_sig_d_not ;
   END LOOP;
end process;

process(clklock_falling_edge_count)
begin
   if(clklock_falling_edge_count >= lock_cyc + 1 and PLL_RST_ipd = '0') then
        SEC_OUT_start <= '1' after clklock_half_period_minus_dly0;
   end if;
end process;

process
begin
   wait until  SEC_OUT_start = '1'; LOOP
      SEC_OUT_sig_3d <= not SEC_OUT_sig_3d;
     wait for clklock_half_period1 * secdiv_p;
      SEC_OUT_sig_3d <= not SEC_OUT_sig_3d ;
     wait for clklock_half_period0 * secdiv_p;
     END LOOP;
end process;

    CLK_OUT_sig_d <= CLK_OUT_sig_d_start and not CLK_OUT_sig_d_not; 

    CLK_OUT_plus_delay <= CLK_OUT_sig_d after tpd when tpd >= 0 ns else
                          CLK_OUT_sig_3d; 

    CLK_OUT <= CLK_OUT_plus_delay and not PLL_RST_ipd;

    PLL_LOCK <= PLL_LOCK_plus and not PLL_RST_ipd when tpd >= 0 ns else
                PLL_LOCK_minus and  not PLL_RST_ipd;

    SEC_OUT_sig_d <=  SEC_OUT_sig_d_start and not SEC_OUT_sig_d_not; 

    SEC_OUT_plus_delay <= SEC_OUT_sig_d after tpd when tpd >= 0 ns else
                          SEC_OUT_sig_3d; 

    SEC_OUT <= SEC_OUT_plus_delay and not PLL_RST_ipd;

end VITAL;

configuration CFG_STDPLLX_VITAL of STDPLLX is 
        for VITAL
        end for; 
end CFG_STDPLLX_VITAL;


----- VITAL model for cell LVDSIN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity LVDSIN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_P_IN_O                      :	VitalDelayType01 := ( 0.00 ns, 0.00 ns);
      tpd_N_IN_O                      :	VitalDelayType01 := ( 0.00 ns, 0.00 ns);
      tipd_N_IN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_P_IN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      N_IN                            :	in    STD_ULOGIC;
      P_IN                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVDSIN : entity is FALSE;
end LVDSIN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of LVDSIN is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL P_IN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (P_IN_ipd, P_IN, tipd_P_IN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (P_IN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(P_IN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (P_IN_ipd'last_event, tpd_P_IN_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell LVDSOUT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity LVDSOUT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I_P_OUT                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_OUT                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I                             :	in    STD_ULOGIC;
      P_OUT                             :	out   STD_ULOGIC;
      N_OUT                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVDSOUT : entity is FALSE;
end LVDSOUT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of LVDSOUT is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(I_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => P_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "P_OUT",
       OutTemp => O_zd,
       Paths => (0 => (I_ipd'last_event, tpd_I_P_OUT, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell LVDSTRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity LVDSTRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_P_OUT                    :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_OE_N_OUT                    :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_I_P_OUT                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_OUT                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_OE                        :	VitalDelayType01 := (0.0 ns, 0.0 ns));

   port(
      I                             :	in    STD_ULOGIC;
      OE                            :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVDSTRI : entity is FALSE;
end LVDSTRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of LVDSTRI is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => I_ipd,
              enable => (NOT OE_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => P_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "P_OUT",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_P_OUT), TRUE),
                 1 => (I_ipd'last_event, VitalExtendToFillDelay(tpd_I_P_OUT), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end LATTICE_ARCH;

----- VITAL model for cell LVDSIO -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity LVDSIO is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_P_IO                      :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_OE_N_IO                      :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_I_P_IO                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_IO                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_P_IO_O                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_N_IO_O                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_OE                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_P_IO                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_N_IO                        :	VitalDelayType01 := (0.0 ns, 0.0 ns));

   port(
      I                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_IO                             :	inout STD_ULOGIC;
      N_IO                             :	inout STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVDSIO : entity is FALSE;
end LVDSIO;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of LVDSIO is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL P_IO_ipd	 : STD_ULOGIC := 'X';
   SIGNAL N_IO_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   VitalWireDelay (P_IO_ipd, P_IO, tipd_P_IO);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd, OE_ipd, P_IO_ipd)


   -- functionality results
--   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
     VARIABLE IO_zd : std_ulogic ;
     VARIABLE O_zd : std_ulogic ;

   -- output glitch detection variables
   VARIABLE IO_GlitchData	: VitalGlitchDataType;
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      IO_zd := VitalBUFIF1 (I_ipd, OE_ipd);
      O_zd := VitalBUF(P_IO_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => P_IO,
       GlitchData => IO_GlitchData,
       OutSignalName => "P_IO",
       OutTemp => IO_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_P_IO), TRUE),
                 1 => (I_ipd'last_event, VitalExtendToFillDelay(tpd_I_P_IO), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (P_IO_ipd'last_event, tpd_P_IO_O, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell BLVDSIN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BLVDSIN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_P_IN_O                      :	VitalDelayType01 := ( 0.00 ns, 0.00 ns);
      tpd_N_IN_O                      :	VitalDelayType01 := ( 0.00 ns, 0.00 ns);
      tipd_N_IN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_P_IN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      N_IN                            :	in    STD_ULOGIC;
      P_IN                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BLVDSIN : entity is FALSE;
end BLVDSIN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of BLVDSIN is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL P_IN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (P_IN_ipd, P_IN, tipd_P_IN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (P_IN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(P_IN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (P_IN_ipd'last_event, tpd_P_IN_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell BLVDSOUT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity BLVDSOUT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I_P_OUT                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_OUT                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I                             :	in    STD_ULOGIC;
      P_OUT                             :	out   STD_ULOGIC;
      N_OUT                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BLVDSOUT : entity is FALSE;
end BLVDSOUT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of BLVDSOUT is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(I_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => P_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "P_OUT",
       OutTemp => O_zd,
       Paths => (0 => (I_ipd'last_event, tpd_I_P_OUT, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell BLVDSTRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BLVDSTRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_P_OUT                    :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_OE_N_OUT                    :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_I_P_OUT                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_OUT                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_OE                        :	VitalDelayType01 := (0.0 ns, 0.0 ns));

   port(
      I                             :	in    STD_ULOGIC;
      OE                            :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BLVDSTRI : entity is FALSE;
end BLVDSTRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of BLVDSTRI is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => I_ipd,
              enable => (NOT OE_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => P_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "P_OUT",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_P_OUT), TRUE),
                 1 => (I_ipd'last_event, VitalExtendToFillDelay(tpd_I_P_OUT), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end LATTICE_ARCH;

----- VITAL model for cell BLVDSIO -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity BLVDSIO is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_P_IO                      :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_OE_N_IO                      :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_I_P_IO                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_IO                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_P_IO_O                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_N_IO_O                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_OE                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_P_IO                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_N_IO                        :	VitalDelayType01 := (0.0 ns, 0.0 ns));

   port(
      I                             :	in    STD_ULOGIC;
      OE                             :	in    STD_ULOGIC;
      P_IO                             :	inout STD_ULOGIC;
      N_IO                             :	inout STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BLVDSIO : entity is FALSE;
end BLVDSIO;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture LATTICE_ARCH of BLVDSIO is
   attribute VITAL_LEVEL1 of LATTICE_ARCH : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL P_IO_ipd	 : STD_ULOGIC := 'X';
   SIGNAL N_IO_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   VitalWireDelay (P_IO_ipd, P_IO, tipd_P_IO);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd, OE_ipd, P_IO_ipd)


   -- functionality results
--   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
     VARIABLE IO_zd : std_ulogic ;
     VARIABLE O_zd : std_ulogic ;

   -- output glitch detection variables
   VARIABLE IO_GlitchData	: VitalGlitchDataType;
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      IO_zd := VitalBUFIF1 (I_ipd, OE_ipd);
      O_zd := VitalBUF(P_IO_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => P_IO,
       GlitchData => IO_GlitchData,
       OutSignalName => "P_IO",
       OutTemp => IO_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_P_IO), TRUE),
                 1 => (I_ipd'last_event, VitalExtendToFillDelay(tpd_I_P_IO), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (P_IO_ipd'last_event, tpd_P_IO_O, TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end LATTICE_ARCH;

----- VITAL model for cell LVPECLIN -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity LVPECLIN is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_P_IN_O                      :	VitalDelayType01 := ( 0.00 ns, 0.00 ns);
      tpd_N_IN_O                      :	VitalDelayType01 := ( 0.00 ns, 0.00 ns);
      tipd_N_IN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_P_IN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      N_IN                            :	in    STD_ULOGIC;
      P_IN                            :	in    STD_ULOGIC;
      O                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVPECLIN : entity is FALSE;
end LVPECLIN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL of LVPECLIN is
   attribute VITAL_LEVEL1 of VITAL : architecture is FALSE;

   SIGNAL P_IN_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (P_IN_ipd, P_IN, tipd_P_IN);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (P_IN_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(P_IN_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => O,
       GlitchData => O_GlitchData,
       OutSignalName => "O",
       OutTemp => O_zd,
       Paths => (0 => (P_IN_ipd'last_event, tpd_P_IN_O, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL;

----- VITAL model for cell LVPECLOUT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity LVPECLOUT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_I_P_OUT                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_OUT                      :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      I                             :	in    STD_ULOGIC;
      P_OUT                             :	out   STD_ULOGIC;
      N_OUT                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVPECLOUT : entity is FALSE;
end LVPECLOUT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL of LVPECLOUT is
   attribute VITAL_LEVEL1 of VITAL : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := TO_X01(I_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => P_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "P_OUT",
       OutTemp => O_zd,
       Paths => (0 => (I_ipd'last_event, tpd_I_P_OUT, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;
end VITAL;

----- VITAL model for cell LVPECLTRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity LVPECLTRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := True;
      MsgOn: Boolean := True;
      tpd_OE_P_OUT                    :	VitalDelayType01Z := (0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns, 0.0 ns);
      tpd_I_P_OUT                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tpd_I_N_OUT                       :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_I                        :	VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_OE                        :	VitalDelayType01 := (0.0 ns, 0.0 ns));

   port(
      I                             :	in    STD_ULOGIC;
      OE                            :	in    STD_ULOGIC;
      P_OUT                          :	out   STD_ULOGIC;
      N_OUT                          :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of LVPECLTRI : entity is FALSE;
end LVPECLTRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;

architecture VITAL of LVPECLTRI is
   attribute VITAL_LEVEL1 of VITAL : architecture is FALSE;

   SIGNAL I_ipd	 : STD_ULOGIC := 'X';
   SIGNAL OE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (I_ipd, I, tipd_I);
   VitalWireDelay (OE_ipd, OE, tipd_OE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (I_ipd, OE_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS O_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE O_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      O_zd := VitalBUFIF0 (data => I_ipd,
              enable => (NOT OE_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => P_OUT,
       GlitchData => O_GlitchData,
       OutSignalName => "P_OUT",
       OutTemp => O_zd,
       Paths => (0 => (OE_ipd'last_event, VitalExtendToFillDelay(tpd_OE_P_OUT), TRUE),
                 1 => (I_ipd'last_event, VitalExtendToFillDelay(tpd_I_P_OUT), TRUE)),
       Mode => VitalInertial,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;
end VITAL;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity AND10 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 Z0 : OUT std_logic);

end AND10;

architecture LATTICE_ARCH of AND10 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND11 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 Z0 : OUT std_logic);

end AND11;

architecture LATTICE_ARCH of AND11 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10)))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND12 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 Z0 : OUT std_logic);

end AND12;

architecture LATTICE_ARCH of AND12 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND13 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 Z0 : OUT std_logic);

end AND13;

architecture LATTICE_ARCH of AND13 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11 AND (A12)))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND14 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 Z0 : OUT std_logic);

end AND14;

architecture LATTICE_ARCH of AND14 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11 AND (A12 AND (A13))))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND15 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 Z0 : OUT std_logic);

end AND15;

architecture LATTICE_ARCH of AND15 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11 AND (A12 AND (A13 AND (A14)))))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND16 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 Z0 : OUT std_logic);

end AND16;

architecture LATTICE_ARCH of AND16 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11 AND (A12 AND (A13 AND (A14 AND (A15))))))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND17 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 A16 : IN std_logic;
		 Z0 : OUT std_logic);

end AND17;

architecture LATTICE_ARCH of AND17 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11 AND (A12 AND (A13 AND (A14 AND (A15 AND (A16)))))))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND18 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 A16 : IN std_logic;
		 A17 : IN std_logic;
		 Z0 : OUT std_logic);

end AND18;

architecture LATTICE_ARCH of AND18 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := A0 AND A1 AND A2 AND A3 AND A4 AND A5 AND A6 AND A7 AND A8 AND A9 AND A10 AND A11 AND A12 AND A13 AND A14 AND A15 AND A16 AND A17;
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND2 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end AND2;

architecture LATTICE_ARCH of AND2 is
begin
		process(A0, A1)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND3 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end AND3;

architecture LATTICE_ARCH of AND3 is
begin
		process(A0, A1, A2)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2)));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND4 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end AND4;

architecture LATTICE_ARCH of AND4 is
begin
		process(A0, A1, A2, A3)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND5 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 Z0 : OUT std_logic);

end AND5;

architecture LATTICE_ARCH of AND5 is
begin
		process(A0, A1, A2, A3, A4)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4)))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND6 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 Z0 : OUT std_logic);

end AND6;

architecture LATTICE_ARCH of AND6 is
begin
		process(A0, A1, A2, A3, A4, A5)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND7 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 Z0 : OUT std_logic);

end AND7;

architecture LATTICE_ARCH of AND7 is
begin
		process(A0, A1, A2, A3, A4, A5, A6)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6)))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND8 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end AND8;

architecture LATTICE_ARCH of AND8 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity AND9 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end AND9;

architecture LATTICE_ARCH of AND9 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8)))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
-------------------------------------------------
--		PRIMITVE BUF UNIT DELAY MODEL		-----
-------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity BUF is

	generic( TDELAY : TIME := 1 ns);

	port (A0 : IN STD_LOGIC;
		  Z0 : OUT STD_LOGIC);
end BUF;


architecture LATTICE_ARCH of BUF is 

begin

	process(A0)

	begin 
			Z0 <= transport A0 after TDELAY;
	end process;

end LATTICE_ARCH;
-------------------------------------------------
--		PRIMITVE FD11 UNIT DELAY MODEL	-----
-------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FD11 is
	generic ( TDELAY : TIME := 1 ns);

 	port( D0, CLK : IN std_logic;
			Q0 : OUT std_logic);

end FD11;

architecture LATTICE_ARCH of FD11 is

begin

	process(D0, CLK)
	variable pQ0 : std_logic;
	variable iQ0 : std_logic;

	begin 

		if CLK'EVENT AND CLK = '1' then
			pQ0 := iQ0;
			if (D0'EVENT) then
				iQ0 := D0'LAST_VALUE;
			elsif NOT(D0'EVENT) then
				iQ0 := D0;
			end if;

			if pQ0 /= iQ0 then
				Q0 <= transport iQ0 after TDELAY;
			else
				Q0 <= transport iQ0;
			end if;

		end if;

	end process;

end LATTICE_ARCH; --// FD11
-------------------------------------------------
--		PRIMITVE FD21 UNIT DELAY MODEL	-----
-------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
entity FD21 is
	generic ( TDELAY : TIME := 1 ns);

 	port( D0, CLK, CD : IN std_logic;
			Q0 : OUT std_logic);


end FD21;


architecture LATTICE_ARCH of FD21 is

begin

	process(D0, CLK, CD)
	variable pQ0 : std_logic;
	variable iQ0 : std_logic;

	begin 

		if CD = '1' then
			if NOT (iQ0 = '0') then
				iQ0 := '0';
				Q0 <= transport iQ0 after TDELAY;
			end if;

		elsif CD = '0' AND CLK'EVENT AND CLK = '1' then
			pQ0 := iQ0;
			if (D0'EVENT) then
				iQ0 := D0'LAST_VALUE;
			elsif NOT(D0'EVENT) then
				iQ0 := D0;
			end if;

			if pQ0 /= iQ0 then
				Q0 <= transport iQ0 after TDELAY;
			else
				Q0 <= transport iQ0;
			end if;

		end if;

	end process;

end LATTICE_ARCH; -- FD21
-------------------------------------------------
--		PRIMITVE INV UNIT DELAY MODEL		-----
-------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity INV is

	generic( TDELAY : TIME := 1 ns);

	port (A0 : IN STD_LOGIC;
		  ZN0 : OUT STD_LOGIC);
end INV;


architecture LATTICE_ARCH of INV is 

begin

	process(A0)

	begin 
			ZN0 <= transport  NOT A0 after TDELAY;
	end process;

end LATTICE_ARCH;
-------------------------------------------------
--		PRIMITVE LXOR2 UNIT DELAY MODEL		-----
-------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity LXOR2 is

	generic( TDELAY : TIME := 1 ns);

	port (A0 : IN STD_LOGIC;
		  A1 : IN STD_LOGIC;
		  Z0 : OUt STD_LOGIC);
end LXOR2;


architecture LATTICE_ARCH of LXOR2 is 

begin

	process(A0, A1)
	variable pZ0 : STD_LOGIC;
	variable iZ0 : STD_LOGIC;

	begin 
		pZ0 := iZ0;
		iZ0 := (A0 XOR A1);
		if pZ0 /= iZ0 then
			Z0 <= transport iZ0 after TDELAY;
		else 
			Z0 <= transport iZ0;
		end if;

	end process;

end LATTICE_ARCH; --// LXOR2
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND10 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND10;

architecture LATTICE_ARCH of NAND10 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND11 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND11;

architecture LATTICE_ARCH of NAND11 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10)))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND12 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND12;

architecture LATTICE_ARCH of NAND12 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11))))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND16 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND16;

architecture LATTICE_ARCH of NAND16 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8 AND (A9 AND (A10 AND (A11 AND (A12 AND (A13 AND (A14 AND (A15))))))))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND2 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND2;

architecture LATTICE_ARCH of NAND2 is
begin
		process(A0, A1)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND3 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND3;

architecture LATTICE_ARCH of NAND3 is
begin
		process(A0, A1, A2)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2)));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND4 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND4;

architecture LATTICE_ARCH of NAND4 is
begin
		process(A0, A1, A2, A3)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND5 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND5;

architecture LATTICE_ARCH of NAND5 is
begin
		process(A0, A1, A2, A3, A4)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4)))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND6 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND6;

architecture LATTICE_ARCH of NAND6 is
begin
		process(A0, A1, A2, A3, A4, A5)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND7 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND7;

architecture LATTICE_ARCH of NAND7 is
begin
		process(A0, A1, A2, A3, A4, A5, A6)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6)))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND8 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND8;

architecture LATTICE_ARCH of NAND8 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NAND9 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end NAND9;

architecture LATTICE_ARCH of NAND9 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 AND (A1 AND (A2 AND (A3 AND (A4 AND (A5 AND (A6 AND (A7 AND (A8)))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR10 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR10;

architecture LATTICE_ARCH of NOR10 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR11 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR11;

architecture LATTICE_ARCH of NOR11 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9 OR (A10)))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR12 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR12;

architecture LATTICE_ARCH of NOR12 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9 OR (A10 OR (A11))))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR16 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR16;

architecture LATTICE_ARCH of NOR16 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9 OR (A10 OR (A11 OR (A12 OR (A13 OR (A14 OR (A15))))))))))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR2 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR2;

architecture LATTICE_ARCH of NOR2 is
begin
		process(A0, A1)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR3 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR3;

architecture LATTICE_ARCH of NOR3 is
begin
		process(A0, A1, A2)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2)));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR4 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR4;

architecture LATTICE_ARCH of NOR4 is
begin
		process(A0, A1, A2, A3)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR5 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR5;

architecture LATTICE_ARCH of NOR5 is
begin
		process(A0, A1, A2, A3, A4)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4)))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR6 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR6;

architecture LATTICE_ARCH of NOR6 is
begin
		process(A0, A1, A2, A3, A4, A5)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR7 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR7;

architecture LATTICE_ARCH of NOR7 is
begin
		process(A0, A1, A2, A3, A4, A5, A6)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6)))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR8 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR8;

architecture LATTICE_ARCH of NOR8 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity NOR9 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end NOR9;

architecture LATTICE_ARCH of NOR9 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8)))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR10 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 Z0 : OUT std_logic);

end OR10;

architecture LATTICE_ARCH of OR10 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR11 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 Z0 : OUT std_logic);

end OR11;

architecture LATTICE_ARCH of OR11 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9 OR (A10)))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR12 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 Z0 : OUT std_logic);

end OR12;

architecture LATTICE_ARCH of OR12 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9 OR (A10 OR (A11))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR16 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 A9 : IN std_logic;
		 A10 : IN std_logic;
		 A11 : IN std_logic;
		 A12 : IN std_logic;
		 A13 : IN std_logic;
		 A14 : IN std_logic;
		 A15 : IN std_logic;
		 Z0 : OUT std_logic);

end OR16;

architecture LATTICE_ARCH of OR16 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8 OR (A9 OR (A10 OR (A11 OR (A12 OR (A13 OR (A14 OR (A15))))))))))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR2 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end OR2;

architecture LATTICE_ARCH of OR2 is
begin
		process(A0, A1)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR3 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end OR3;

architecture LATTICE_ARCH of OR3 is
begin
		process(A0, A1, A2)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2)));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR4 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end OR4;

architecture LATTICE_ARCH of OR4 is
begin
		process(A0, A1, A2, A3)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR5 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 Z0 : OUT std_logic);

end OR5;

architecture LATTICE_ARCH of OR5 is
begin
		process(A0, A1, A2, A3, A4)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4)))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR6 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 Z0 : OUT std_logic);

end OR6;

architecture LATTICE_ARCH of OR6 is
begin
		process(A0, A1, A2, A3, A4, A5)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR7 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 Z0 : OUT std_logic);

end OR7;

architecture LATTICE_ARCH of OR7 is
begin
		process(A0, A1, A2, A3, A4, A5, A6)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6)))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR8 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end OR8;

architecture LATTICE_ARCH of OR8 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity OR9 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end OR9;

architecture LATTICE_ARCH of OR9 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 OR (A1 OR (A2 OR (A3 OR (A4 OR (A5 OR (A6 OR (A7 OR (A8)))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;


entity PW is

	port( PULSE : IN std_logic);

end PW;

architecture LATTICE_ARCH of PW is

begin

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;


entity SHFE is

	port( REF : IN std_logic;
		DATA : IN std_logic);

end SHFE;

architecture LATTICE_ARCH of SHFE is

begin

end LATTICE_ARCH; -- SHFE

-------------------------------------------------
--		PRIMITVE XBIDI UNIT DELAY MODEL	-----
-------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XBIDI1 is
	
	generic ( TDELAY : TIME := 1 ns);
	port ( A0 : IN std_logic;
		   OE : IN std_logic;
		   Z0 : OUT std_logic;
		   XB0 : INOUT std_logic);

end XBIDI1;

architecture LATTICE_ARCH of XBIDI1 is

begin

	process(A0, OE, XB0)
	variable pZ0 : std_logic;
	variable iZ0 : std_logic;

	begin

	pZ0 := iZ0;
	if OE = '1' then
		iZ0 := A0;
		if pZ0 /= iZ0 then
			XB0 <= transport iZ0 after TDELAY;
			Z0 <= transport iZ0 after TDELAY;
		else 
			XB0 <= transport iZ0 ;
			Z0 <= transport iZ0 ;
		end if;
	elsif OE = '0' then
		iZ0 := 'Z';
		if pZ0 /= iZ0 then
			XB0 <= transport iZ0 after TDELAY;
			Z0 <= transport XB0 after TDELAY;
		else 
			XB0 <= transport iZ0 ;
			Z0 <= transport XB0 ;
		end if;
	end if;

	end process;

end LATTICE_ARCH;

-------------------------------------------------
--		PRIMITVE XDFF1 UNIT DELAY MODEL	-----
-------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity XDFF1 is
	generic ( TDELAY : TIME := 1 ns);

 	port( D0, CLK : IN std_logic;
			Q0 : OUT std_logic);
end XDFF1;

architecture LATTICE_ARCH of XDFF1 is

begin

	process(D0, CLK)
	variable pQ0 : std_logic;
	variable iQ0 : std_logic;

	begin 

		if CLK'EVENT AND CLK = '1' then
			pQ0 := iQ0;
			if (D0'EVENT) then
				iQ0 := D0'LAST_VALUE;
			elsif NOT(D0'EVENT) then
				iQ0 := D0;
			end if;

			if pQ0 /= iQ0 then
				Q0 <= transport iQ0 after TDELAY;
			else
				Q0 <= transport iQ0;
			end if;

		end if;


	end process;

end LATTICE_ARCH;-- XDFF1
-------------------------------------------------
--		PRIMITVE XDL1 UNIT DELAY MODEL	-----
-------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XDL1 is
	
		generic ( TDELAY : TIME := 1 ns);
		port ( D0 : IN std_logic;
				G : IN std_logic;
			   Q0 : OUT std_logic);
end XDL1;

architecture LATTICE_ARCH of XDL1 is

begin

	process(D0, G)

	variable pQ0 : std_logic;
	variable iQ0 : std_logic;
				
	begin

	pQ0 := iQ0;

	if G = '1' then

		iQ0 := D0;
		if pQ0 /= iQ0 then
			Q0 <= transport iQ0 after TDELAY;
		else 
			Q0 <= transport iQ0;
		end if;

	end if;
		
	end process;

end LATTICE_ARCH;
-------------------------------------------------
--		PRIMITVE XINPUT UNIT DELAY MODEL	-----
-------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity XINPUT is

	generic( TDELAY : TIME := 1 ns);

	port( XI0 : IN  STD_LOGIC;
		  Z0  : OUT STD_LOGIC);

end XINPUT;


architecture LATTICE_ARCH of XINPUT is

begin

	process(XI0)

	begin 
			Z0 <= transport XI0 after TDELAY;
	end process;

--	component BUF
--		port( A0 : IN std_logic;
--			  Z0 : OUT std_logic);
--end component;

--begin
--	UQXIN : BUF
--		port map (Z0 => Z0, A0 => XI0);

end LATTICE_ARCH; -- XINPUT
-------------------------------------------------
--		PRIMITVE XINV UNIT DELAY MODEL		-----
-------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity XINV is

	generic( TDELAY : TIME := 1 ns);

	port (A0 : IN STD_LOGIC;
		  ZN0 : OUT STD_LOGIC);
end XINV;


architecture LATTICE_ARCH of XINV is 

begin

	process(A0)

	begin 
			ZN0 <= transport  NOT A0 after TDELAY;
	end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XNOR2 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 ZN0 : OUT std_logic);

end XNOR2;

architecture LATTICE_ARCH of XNOR2 is
begin
		process(A0, A1)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT( A0 XOR (A1));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XNOR3 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 ZN0 : OUT std_logic);

end XNOR3;

architecture LATTICE_ARCH of XNOR3 is
begin
		process(A0, A1, A2)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT( A0 XOR (A1 XOR (A2)));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XNOR4 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 ZN0 : OUT std_logic);

end XNOR4;

architecture LATTICE_ARCH of XNOR4 is
begin
		process(A0, A1, A2, A3)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT( A0 XOR (A1 XOR (A2 XOR (A3))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XNOR7 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 ZN0 : OUT std_logic);

end XNOR7;

architecture LATTICE_ARCH of XNOR7 is
begin
		process(A0, A1, A2, A3, A4, A5, A6)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT( A0 XOR (A1 XOR (A2 XOR (A3 XOR (A4 XOR (A5 XOR (A6)))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XNOR8 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 ZN0 : OUT std_logic);

end XNOR8;

architecture LATTICE_ARCH of XNOR8 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT( A0 XOR (A1 XOR (A2 XOR (A3 XOR (A4 XOR (A5 XOR (A6 XOR (A7))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XNOR9 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 ZN0 : OUT std_logic);

end XNOR9;

architecture LATTICE_ARCH of XNOR9 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := NOT( A0 XOR (A1 XOR (A2 XOR (A3 XOR (A4 XOR (A5 XOR (A6 XOR (A7 XOR (A8)))))))));
			if pZ0 /= iZ0 then
				ZN0 <= transport iZ0 after TDELAY;
			else
				ZN0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XOR2 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 Z0 : OUT std_logic);

end XOR2;

architecture LATTICE_ARCH of XOR2 is
begin
		process(A0, A1)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 XOR (A1));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XOR3 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 Z0 : OUT std_logic);

end XOR3;

architecture LATTICE_ARCH of XOR3 is
begin
		process(A0, A1, A2)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 XOR (A1 XOR (A2)));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XOR4 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 Z0 : OUT std_logic);

end XOR4;

architecture LATTICE_ARCH of XOR4 is
begin
		process(A0, A1, A2, A3)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 XOR (A1 XOR (A2 XOR (A3))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XOR8 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 Z0 : OUT std_logic);

end XOR8;

architecture LATTICE_ARCH of XOR8 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 XOR (A1 XOR (A2 XOR (A3 XOR (A4 XOR (A5 XOR (A6 XOR (A7))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


entity XOR9 is
	generic ( TDELAY : TIME := 1 ns);
	port(A0 : IN std_logic;
		 A1 : IN std_logic;
		 A2 : IN std_logic;
		 A3 : IN std_logic;
		 A4 : IN std_logic;
		 A5 : IN std_logic;
		 A6 : IN std_logic;
		 A7 : IN std_logic;
		 A8 : IN std_logic;
		 Z0 : OUT std_logic);

end XOR9;

architecture LATTICE_ARCH of XOR9 is
begin
		process(A0, A1, A2, A3, A4, A5, A6, A7, A8)
		variable pZ0 : std_logic;
		variable iZ0 : std_logic;

		 begin
			pZ0 := iZ0;
			iZ0 := (A0 XOR (A1 XOR (A2 XOR (A3 XOR (A4 XOR (A5 XOR (A6 XOR (A7 XOR (A8)))))))));
			if pZ0 /= iZ0 then
				Z0 <= transport iZ0 after TDELAY;
			else
				Z0 <= transport iZ0;
			end if;
		end process;

end LATTICE_ARCH;
-------------------------------------------------
--		PRIMITVE XOUTPUT UNIT DELAY MODEL	-----
-------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity XOUTPUT is

	generic( TDELAY : TIME := 1 ns);

	port( A0 : IN  STD_LOGIC;
		  XO0  : OUT STD_LOGIC);

end XOUTPUT;


architecture LATTICE_ARCH of XOUTPUT is

begin

	process(A0)

	begin 
			XO0 <= transport A0 after TDELAY;
	end process;

--	component BUF
--		port( A0 : IN std_logic;
--			  Z0 : OUT std_logic);

--end component;

--begin

--	UQXOUT : BUF
--		port map (Z0 => XO0, A0 => A0);

end LATTICE_ARCH; -- XOUTPUT


-------------------------------------------------
--		PRIMITVE XTRI1 UNIT DELAY MODEL	-----
-------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
entity XTRI1 is

	generic ( TDELAY : TIME := 1 ns);

	port( A0 : IN  std_logic;
		  OE : IN  std_logic;
		  XO0 : OUT  std_logic);

end XTRI1;

architecture LATTICE_ARCH of XTRI1 is

begin

	process(A0, OE)

	variable pXO0 : std_logic;
	variable iXO0 : std_logic;

	begin

		pXO0 := iXO0;
		if OE'EVENT AND OE = '1' then
			iXO0 := A0;
			if pXO0 /= iXO0 then
				XO0 <=  transport iXO0 after TDELAY;
			else
				XO0 <= transport iXO0;
			end if;

		elsif OE'EVENT AND OE = '0' then
			iXO0 := 'Z';
			if pXO0 /= iXO0 then
				XO0 <=  transport iXO0 after TDELAY;
			else
				XO0 <= transport iXO0;
			end if;

		elsif A0'EVENT  AND OE = '1' then
			iXO0 := A0;
			if pXO0 /= iXO0 then
				XO0 <=  transport iXO0 after TDELAY;
			else 
				XO0 <= transport iXO0;
			end if;   

		end if;
	end process;

end LATTICE_ARCH; -- XTRI1
--*****************************************************--
--   The following primitives are built for 8K device  --
--   while unit delay is used                          --
--*****************************************************--

Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FD11E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, EN : IN std_logic;
	       Q0 : OUT std_logic);
end FD11E;

architecture LATTICE_ARCH of FD11E is

signal iD0 : std_logic;

begin

  process(D0, CLK, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin

    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);

    if CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;

       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FD21E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end FD21E;

architecture LATTICE_ARCH of FD21E is

signal iD0 : std_logic;

begin

  process(D0, CLK, CD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);

    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;

       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FDC1 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end FDC1;

architecture LATTICE_ARCH of FDC1 is

begin

  process(D0, CLK, SD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    
    if SD = '1' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (D0'EVENT) then
	iQ0 := D0'last_value;
       elsif NOT(D0'EVENT) then
	iQ0 := D0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FDC1E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, SD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end FDC1E;

architecture LATTICE_ARCH of FDC1E is

signal iD0 : std_logic;

begin

  process(D0, CLK, SD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);
    
    if SD = '1' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FDE1 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD, SD : IN std_logic;
	           Q0 : OUT std_logic);
end FDE1;

architecture LATTICE_ARCH of FDE1 is

begin

  process(D0, CLK, CD, SD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    
    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (D0'EVENT) then
	iQ0 := D0'last_value;
       elsif NOT(D0'EVENT) then
	iQ0 := D0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FDE1E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD, SD, EN : IN std_logic;
	               Q0 : OUT std_logic);
end FDE1E;

architecture LATTICE_ARCH of FDE1E is

signal iD0 : std_logic;

begin

  process(D0, CLK, CD, SD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);
    
    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FTI21 is
  generic (TDELAY : TIME := 1 ns);
  port (T0, CLK, CD : IN std_logic;
                 Q0 : OUT std_logic);
end FTI21;

architecture LATTICE_ARCH of FTI21 is
begin

  process(T0, CLK, CD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin

    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND CLK'EVENT AND CLK='1' then
       pQ0 := iQ0;
       if (T0'EVENT) then
	iQ0 := T0'last_value XOR iQ0;
       elsif NOT(T0'EVENT) then
	iQ0 := T0 XOR iQ0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;

     end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FTI21E is
  generic (TDELAY : TIME := 1 ns);
  port (T0, CLK, CD, EN : IN std_logic;
                     Q0 : OUT std_logic);
end FTI21E;

architecture LATTICE_ARCH of FTI21E is

signal iT0 : std_logic;

begin

  process(T0, CLK, CD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iT0 <= T0 AND EN;

    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND CLK'EVENT AND CLK='1' then
       pQ0 := iQ0;
       if (iT0'EVENT) then
	iQ0 := iT0'last_value XOR iQ0;
       else
	iQ0 := iT0 XOR iQ0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;

    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FTI31 is
  generic (TDELAY : TIME := 1 nS);
  port (T0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end FTI31;

architecture LATTICE_ARCH of FTI31 is
begin

  process(T0, CLK, SD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin

    if SD = '1' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (T0'EVENT) then
	iQ0 := T0'last_value XOR iQ0;
       elsif NOT(T0'EVENT) then
	iQ0 := T0 XOR iQ0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;

     end if;
   end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FTI31E is
  generic (TDELAY : TIME := 1 ns);
  port (T0, CLK, SD, EN : IN std_logic;
		 Q0 : OUT std_logic);
end FTI31E;

architecture LATTICE_ARCH of FTI31E is

signal iT0 : std_logic;

begin

  process(T0, CLK, SD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iT0 <= T0 AND EN;

    if SD = '1' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (iT0'EVENT) then
	iQ0 := iT0'last_value XOR iQ0;
       else
	iQ0 := iT0 XOR iQ0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;

     end if;
   end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FTI41 is
  generic (TDELAY : TIME := 1 ns);
  port (T0, CLK, SD, CD : IN std_logic;
		 Q0 : OUT std_logic);
end FTI41;

architecture LATTICE_ARCH of FTI41 is
begin

  process(T0, CLK, SD, CD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin

    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (T0'EVENT) then
	iQ0 := T0'last_value XOR iQ0;
       elsif NOT(T0'EVENT) then
	iQ0 := T0 XOR iQ0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;

     end if;
   end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity FTI41E is
  generic (TDELAY : TIME := 1 ns);
  port (T0, CLK, CD, SD, EN : IN std_logic;
		     Q0 : OUT std_logic);
end FTI41E;

architecture LATTICE_ARCH of FTI41E is

signal iT0 : std_logic;

begin

  process(T0, CLK, SD, CD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iT0 <= T0 AND EN;

    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (iT0'EVENT) then
	iQ0 := iT0'last_value XOR iQ0;
       else
          iQ0 := iT0 XOR iQ0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;

    end if;
  end process;

end LATTICE_ARCH;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

entity IT11 is
  generic (TDELAY : TIME := 1 ns);
  port(A0, OE : IN std_logic;
	 O0 : OUT  std_logic);
end IT11;
       
architecture LATTICE_ARCH of IT11 is
begin

  process(A0, OE)
  variable pO0 : std_logic;
  variable iO0 : std_logic;
  begin
    pO0 := iO0;

    if OE'EVENT AND OE = '1' then
      iO0 := A0;
      if pO0 /= iO0 then
        O0 <=  transport iO0 after TDELAY;
      else
        O0 <= transport iO0;
      end if;

    elsif OE'EVENT AND OE = '0' then
      iO0 := 'Z';
      if pO0 /= iO0 then
        O0 <=  transport iO0 after TDELAY;
      else
        O0 <= transport iO0;
      end if;

    elsif A0'EVENT  AND OE = '1' then
      iO0 := A0;
      if pO0 /= iO0 then
        O0 <=  transport iO0 after TDELAY;
      else
        O0 <= transport iO0;
      end if;

    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity LDI11 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G : IN std_logic;
           Q0 : OUT std_logic);
end LDI11;

architecture LATTICE_ARCH of LDI11 is

begin

  process(D0, G)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    pQ0 := iQ0;

    if G = '1' then
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity LDI21 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G, CD : IN std_logic;
	     Q0 : OUT std_logic);
end LDI21;

architecture LATTICE_ARCH of LDI21 is

begin

  process(D0, G, CD)
  variable iQ0 : std_logic;
  variable pQ0 : std_logic;
  begin

    if CD = '1' then
       if NOT(iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;
    
    elsif CD = '0' AND G = '1' then
       pQ0 := iQ0;
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity LDI31 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G, SD : IN std_logic;
	     Q0 : OUT std_logic);
end LDI31;

architecture LATTICE_ARCH of LDI31 is

begin

  process(D0, G, SD)
  variable iQ0 : std_logic;
  variable pQ0 : std_logic;
  begin

    if SD = '1' then
       if NOT(iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;
    
    elsif SD = '0' AND G = '1' then
       pQ0 := iQ0;
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity LDI41 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G, CD, SD : IN std_logic;
	         Q0 : OUT std_logic);
end LDI41;

architecture LATTICE_ARCH of LDI41 is

begin

  process(D0, G, SD, CD)
  variable iQ0 : std_logic;
  variable pQ0 : std_logic;
  begin

    if CD = '1' then
       if NOT(iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT(iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;
    
    elsif CD = '0' AND SD = '0' AND G = '1' then
       pQ0 := iQ0;
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF1E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, EN : IN std_logic;
	       Q0 : OUT std_logic);
end XDFF1E;

architecture LATTICE_ARCH of XDFF1E is

signal iD0 : std_logic;

begin

  process(D0, CLK, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin

    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);

    if CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;

       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF2 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD : IN std_logic;
	       Q0 : OUT std_logic);
end XDFF2;

architecture LATTICE_ARCH of XDFF2 is

begin

  process(D0, CLK, CD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    if CD = '1' then
       if NOT (iQ0 = '0') then
          iQ0 := '0';
          Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (D0'EVENT) then
          iQ0 := D0'last_value;
       elsif NOT(D0'EVENT) then
          iQ0 := D0;
       end if;

       if pQ0 /= iQ0 then
          Q0 <= transport iQ0 after TDELAY;
       else
          Q0 <= transport iQ0;
       end if;

    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF2E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end XDFF2E;

architecture LATTICE_ARCH of XDFF2E is

  signal iD0 : std_logic;

begin

  process(D0, CLK, CD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);

    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;

       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF3 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, SD : IN std_logic;
	       Q0 : OUT std_logic);
end XDFF3;

architecture LATTICE_ARCH of XDFF3 is

begin

  process(D0, CLK, SD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    
    if SD = '1' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (D0'EVENT) then
	iQ0 := D0'last_value;
       elsif NOT(D0'EVENT) then
	iQ0 := D0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF3E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, SD, EN : IN std_logic;
	           Q0 : OUT std_logic);
end XDFF3E;

architecture LATTICE_ARCH of XDFF3E is

  signal iD0 : std_logic;

begin

  process(D0, CLK, SD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);
    
    if SD = '1' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF4 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD, SD : IN std_logic;
	           Q0 : OUT std_logic);
end XDFF4;

architecture LATTICE_ARCH of XDFF4 is

begin

  process(D0, CLK, CD, SD)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    
    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (D0'EVENT) then
	iQ0 := D0'last_value;
       elsif NOT(D0'EVENT) then
	iQ0 := D0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDFF4E is
  generic (TDELAY : TIME := 1 ns);
  port (D0, CLK, CD, SD, EN : IN std_logic;
	               Q0 : OUT std_logic);
end XDFF4E;

architecture LATTICE_ARCH of XDFF4E is

  signal iD0 : std_logic;

begin

  process(D0, CLK, CD, SD, EN)
  variable pQ0 : std_logic;
  variable iQ0 : std_logic;
  begin
    iD0 <= (D0 AND EN) OR (iQ0 AND NOT EN);
    
    if CD = '1' then
       if NOT (iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT (iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif CD = '0' AND SD = '0' AND CLK'EVENT AND CLK = '1' then
       pQ0 := iQ0;
       if (iD0'EVENT) then
	iQ0 := iD0'last_value;
       elsif NOT(iD0'EVENT) then
	iQ0 := iD0;
       end if;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;

  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDL2 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G, CD : IN std_logic;
	     Q0 : OUT std_logic);
end XDL2;

architecture LATTICE_ARCH of XDL2 is

begin

  process(D0, G, CD)
  variable iQ0 : std_logic;
  variable pQ0 : std_logic;
  begin

    if CD = '1' then
       if NOT(iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;
    
    elsif CD = '0' AND G = '1' then
       pQ0 := iQ0;
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDL3 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G, SD : IN std_logic;
	     Q0 : OUT std_logic);
end XDL3;

architecture LATTICE_ARCH of XDL3 is

begin

  process(D0, G, SD)
  variable iQ0 : std_logic;
  variable pQ0 : std_logic;
  begin

    if SD = '1' then
       if NOT(iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;
    
    elsif SD = '0' AND G = '1' then
       pQ0 := iQ0;
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;
Library IEEE;
Use IEEE.STD_LOGIC_1164.all;

entity XDL4 is
  generic (TDELAY : TIME := 1 ns);
  port (D0, G, CD, SD : IN std_logic;
	         Q0 : OUT std_logic);
end XDL4;

architecture LATTICE_ARCH of XDL4 is

begin

  process(D0, G, SD, CD)
  variable iQ0 : std_logic;
  variable pQ0 : std_logic;
  begin

    if CD = '1' then
       if NOT(iQ0 = '0') then
	iQ0 := '0';
	Q0 <= transport iQ0 after TDELAY;
       end if;

    elsif SD = '1' AND CD = '0' then
       if NOT(iQ0 = '1') then
	iQ0 := '1';
	Q0 <= transport iQ0 after TDELAY;
       end if;
    
    elsif CD = '0' AND SD = '0' AND G = '1' then
       pQ0 := iQ0;
       iQ0 := D0;

       if pQ0 /= iQ0 then
	Q0 <= transport iQ0 after TDELAY;
       else
	Q0 <= transport iQ0;
       end if;
    end if;
  end process;

end LATTICE_ARCH;

--*********************************************************
--	This file contains the VHDL source of the macros
--	of the lattice library.
--*********************************************************

-- VHDL netlist for ADDF1
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDF1 IS 
    PORT (
        A0 : IN std_logic;
        B0 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDF1;


ARCHITECTURE lattice_arch OF ADDF1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => CI);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => B0, A1 => UQVN_N1);
UQVB_B3 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N3, A1 => UQVN_N2);
UQVB_B4 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N4);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => B0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => CI);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => CI, A1 => B0);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => CI, A1 => A0);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => B0, A1 => A0);
UQVB_B10 : OR3
	PORT MAP (Z0 => CO, A0 => UQVN_N5, A1 => UQVN_N6, A2 => UQVN_N7);
END lattice_arch;
-- VHDL netlist for ADDF16A
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDF16A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B10 : IN std_logic;
        B11 : IN std_logic;
        B12 : IN std_logic;
        B13 : IN std_logic;
        B14 : IN std_logic;
        B15 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        B8 : IN std_logic;
        B9 : IN std_logic;
        CI : IN std_logic;
        CO : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z10 : OUT std_logic;
        Z11 : OUT std_logic;
        Z12 : OUT std_logic;
        Z13 : OUT std_logic;
        Z14 : OUT std_logic;
        Z15 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        Z8 : OUT std_logic;
        Z9 : OUT std_logic
    );
END ADDF16A;


ARCHITECTURE lattice_arch OF ADDF16A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 UQVN_N113, UQVN_N114, UQVN_N115, UQVN_N116,
	 UQVN_N117, UQVN_N118, UQVN_N119, UQVN_N120,
	 UQVN_N121, UQVN_N122, UQVN_N123, UQVN_N124,
	 UQVN_N125, UQVN_N126, UQVN_N127, UQVN_N128,
	 UQVN_N129, UQVN_N130, UQVN_N131, UQVN_N132,
	 UQVN_N133, UQVN_N134, UQVN_N135, UQVN_N136,
	 UQVN_N137, UQVN_N138, UQVN_N139, UQVN_N140,
	 UQVN_N141, UQVN_N142, UQVN_N143, UQVN_N144,
	 UQVN_N145, UQVN_N146, UQVN_N147, UQVN_N148,
	 UQVN_N149, UQVN_N150, UQVN_N151, UQVN_N152,
	 UQVN_N153, UQVN_N154, UQVN_N155, UQVN_N156,
	 UQVN_N157, UQVN_N158, UQVN_N159, UQVN_N160,
	 UQVN_N161, UQVN_N162, UQVN_N163, UQVN_N164,
	 UQVN_N165, UQVN_N166, UQVN_N167, UQVN_N168,
	 UQVN_N169, UQVN_N170, UQVN_N171, UQVN_N172,
	 UQVN_N173, UQVN_N174, UQVN_N175, UQVN_N176,
	 UQVN_N177, UQVN_N178, UQVN_N179, UQVN_N180,
	 UQVN_N181, UQVN_N182, UQVN_N183, UQVN_N184,
	 UQVN_N185, UQVN_N186, UQVN_N187, UQVN_N188,
	 UQVN_N189, UQVN_N190, UQVN_N191, UQVN_N192,
	 UQVN_N193, UQVN_N194, UQVN_N195, UQVN_N196,
	 UQVN_N197, UQVN_N198, UQVN_N199, UQVN_N200,
	 UQVN_N201, UQVN_N202, UQVN_N203, UQVN_N204,
	 UQVN_N205, UQVN_N206, UQVN_N207, UQVN_N208,
	 UQVN_N209, UQVN_N210, UQVN_N211, UQVN_N212,
	 UQVN_N213, UQVN_N214, UQVN_N215, UQVN_N216,
	 UQVN_N217, UQVN_N218, UQVN_N219, UQVN_N220,
	 UQVN_N221, UQVN_N222, UQVN_N223, UQVN_N224,
	 UQVN_N225, UQVN_N226, UQVN_N227, UQVN_N228,
	 UQVN_N229, UQVN_N230, UQVN_N231, UQVN_N232,
	 UQVN_N233, UQVN_N234, UQVN_N235, UQVN_N236,
	 UQVN_N237, UQVN_N238, UQVN_N239, G012,
	 G1214, G345, G678, G911,
	 P012, P1214, P345, P678,
	 P911 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => P345, A1 => UQVN_N239);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N235, A0 => G345, A1 => UQVN_N1);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N236, A0 => G678, A1 => UQVN_N2, A2 => UQVN_N3);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => P678, A1 => P345, A2 => UQVN_N239);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => P678, A1 => G345);
UQVB_B6 : OR4
	PORT MAP (Z0 => UQVN_N237, A0 => G911, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => UQVN_N6);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => P911, A1 => G678);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => P911, A1 => P678, A2 => G345);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => P911, A1 => P678, A2 => P345, 
	A3 => UQVN_N239);
UQVB_B10 : OR5
	PORT MAP (Z0 => UQVN_N238, A0 => G1214, A1 => UQVN_N7, A2 => UQVN_N8, 
	A3 => UQVN_N9, A4 => UQVN_N10);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => P1214, A1 => G911);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => P1214, A1 => P911, A2 => G678);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => G345);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => P345, A4 => UQVN_N239);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => P012, A1 => CI);
UQVB_B16 : OR2
	PORT MAP (Z0 => UQVN_N239, A0 => G012, A1 => UQVN_N11);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => CI);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => B1);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => B2);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => A0);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N51, A1 => CI);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => B0, A1 => UQVN_N54);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N12, A1 => UQVN_N13);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N14);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N48, A1 => B1, A2 => UQVN_N51);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N52, A1 => B0, A2 => CI);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => A0, A1 => UQVN_N52, A2 => CI);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => B1, A1 => UQVN_N51, A2 => UQVN_N54);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N48, A1 => B1, A2 => UQVN_N54);
UQVB_B30 : OR6
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N15, 
	A3 => UQVN_N16, A4 => UQVN_N20, A5 => UQVN_N19);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N21);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => A0, A1 => UQVN_N52, A2 => B0);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => A0, A1 => A1, A2 => A2, 
	A3 => B0);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => A1, A1 => A2, A2 => B1);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => A0, A1 => A2, A2 => B0, 
	A3 => B1);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => A2, A1 => B2);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B2);
UQVB_B38 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => A1, A1 => B1, A2 => B2);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A0, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B40 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N22, A4 => UQVN_N26, A5 => UQVN_N27, A6 => UQVN_N28);
UQVB_B41 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N48, A1 => UQVN_N51);
UQVB_B42 : AND2
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N49, A1 => UQVN_N52);
UQVB_B43 : AND2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N50, A1 => UQVN_N53);
UQVB_B44 : NOR3
	PORT MAP (ZN0 => P012, A0 => UQVN_N31, A1 => UQVN_N29, A2 => UQVN_N30);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => B0);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => A1);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => A2);
UQVB_B48 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N45);
UQVB_B49 : AND4
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N51, A1 => UQVN_N52, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B50 : AND4
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N48, A1 => UQVN_N52, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N49, A1 => UQVN_N51, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B52 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N48, A1 => UQVN_N49, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B53 : AND4
	PORT MAP (Z0 => UQVN_N41, A0 => B0, A1 => B1, A2 => UQVN_N53, 
	A3 => CI);
UQVB_B54 : AND4
	PORT MAP (Z0 => UQVN_N40, A0 => A0, A1 => B1, A2 => UQVN_N53, 
	A3 => CI);
UQVB_B55 : AND4
	PORT MAP (Z0 => UQVN_N39, A0 => A1, A1 => B0, A2 => UQVN_N53, 
	A3 => CI);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => A0, A1 => A1, A2 => UQVN_N53, 
	A3 => CI);
UQVB_B57 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => A0, A1 => B0, A2 => B1, 
	A3 => UQVN_N53);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N36, A0 => A1, A1 => B1, A2 => UQVN_N53);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => A0, A1 => A1, A2 => B0, 
	A3 => UQVN_N53);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N48, A1 => UQVN_N51, A2 => UQVN_N52, 
	A3 => B2);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N49, A1 => UQVN_N52, A2 => B2);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N48, A1 => UQVN_N49, A2 => UQVN_N51, 
	A3 => B2);
UQVB_B63 : OR12
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N43, A1 => UQVN_N42, A2 => UQVN_N41, 
	A3 => UQVN_N40, A4 => UQVN_N39, A5 => UQVN_N38, A6 => UQVN_N37, 
	A7 => UQVN_N36, A8 => UQVN_N35, A9 => UQVN_N34, A10 => UQVN_N33, 
	A11 => UQVN_N32);
UQVB_B64 : OR3
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N44, A1 => UQVN_N46, A2 => UQVN_N47);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N97, A0 => UQVN_N239);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N95, A0 => B4);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N96, A0 => B5);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N91, A0 => A3);
UQVB_B69 : AND2
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N94, A1 => UQVN_N239);
UQVB_B70 : AND2
	PORT MAP (Z0 => UQVN_N56, A0 => B3, A1 => UQVN_N97);
UQVB_B71 : OR2
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N55, A1 => UQVN_N56);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N57);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N91, A1 => B4, A2 => UQVN_N94);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N95, A1 => B3, A2 => UQVN_N239);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => A3, A1 => UQVN_N95, A2 => UQVN_N239);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N60, A0 => B4, A1 => UQVN_N94, A2 => UQVN_N97);
UQVB_B77 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N91, A1 => B4, A2 => UQVN_N97);
UQVB_B78 : OR6
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N61, A1 => UQVN_N60, A2 => UQVN_N58, 
	A3 => UQVN_N59, A4 => UQVN_N63, A5 => UQVN_N62);
UQVB_B79 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N64);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => A3, A1 => UQVN_N95, A2 => B3);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N68, A0 => A3, A1 => A4, A2 => A5, 
	A3 => B3);
UQVB_B82 : AND3
	PORT MAP (Z0 => UQVN_N67, A0 => A4, A1 => A5, A2 => B4);
UQVB_B83 : AND4
	PORT MAP (Z0 => UQVN_N66, A0 => A3, A1 => A5, A2 => B3, 
	A3 => B4);
UQVB_B84 : AND2
	PORT MAP (Z0 => UQVN_N65, A0 => A5, A1 => B5);
UQVB_B85 : AND4
	PORT MAP (Z0 => UQVN_N69, A0 => A3, A1 => A4, A2 => B3, 
	A3 => B5);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N70, A0 => A4, A1 => B4, A2 => B5);
UQVB_B87 : AND4
	PORT MAP (Z0 => UQVN_N71, A0 => A3, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B88 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N68, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => UQVN_N65, A4 => UQVN_N69, A5 => UQVN_N70, A6 => UQVN_N71);
UQVB_B89 : AND2
	PORT MAP (Z0 => UQVN_N74, A0 => UQVN_N91, A1 => UQVN_N94);
UQVB_B90 : AND2
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N92, A1 => UQVN_N95);
UQVB_B91 : AND2
	PORT MAP (Z0 => UQVN_N73, A0 => UQVN_N93, A1 => UQVN_N96);
UQVB_B92 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N74, A1 => UQVN_N72, A2 => UQVN_N73);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N94, A0 => B3);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N92, A0 => A4);
UQVB_B95 : INV
	PORT MAP (ZN0 => UQVN_N93, A0 => A5);
UQVB_B96 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N88);
UQVB_B97 : AND4
	PORT MAP (Z0 => UQVN_N87, A0 => UQVN_N94, A1 => UQVN_N95, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B98 : AND4
	PORT MAP (Z0 => UQVN_N89, A0 => UQVN_N91, A1 => UQVN_N95, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B99 : AND4
	PORT MAP (Z0 => UQVN_N86, A0 => UQVN_N92, A1 => UQVN_N94, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B100 : AND4
	PORT MAP (Z0 => UQVN_N85, A0 => UQVN_N91, A1 => UQVN_N92, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B101 : AND4
	PORT MAP (Z0 => UQVN_N84, A0 => B3, A1 => B4, A2 => UQVN_N96, 
	A3 => UQVN_N239);
UQVB_B102 : AND4
	PORT MAP (Z0 => UQVN_N83, A0 => A3, A1 => B4, A2 => UQVN_N96, 
	A3 => UQVN_N239);
UQVB_B103 : AND4
	PORT MAP (Z0 => UQVN_N82, A0 => A4, A1 => B3, A2 => UQVN_N96, 
	A3 => UQVN_N239);
UQVB_B104 : AND4
	PORT MAP (Z0 => UQVN_N81, A0 => A3, A1 => A4, A2 => UQVN_N96, 
	A3 => UQVN_N239);
UQVB_B105 : AND4
	PORT MAP (Z0 => UQVN_N80, A0 => A3, A1 => B3, A2 => B4, 
	A3 => UQVN_N96);
UQVB_B106 : AND3
	PORT MAP (Z0 => UQVN_N79, A0 => A4, A1 => B4, A2 => UQVN_N96);
UQVB_B107 : AND4
	PORT MAP (Z0 => UQVN_N78, A0 => A3, A1 => A4, A2 => B3, 
	A3 => UQVN_N96);
UQVB_B108 : AND4
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N91, A1 => UQVN_N94, A2 => UQVN_N95, 
	A3 => B5);
UQVB_B109 : AND3
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N92, A1 => UQVN_N95, A2 => B5);
UQVB_B110 : AND4
	PORT MAP (Z0 => UQVN_N75, A0 => UQVN_N91, A1 => UQVN_N92, A2 => UQVN_N94, 
	A3 => B5);
UQVB_B111 : OR12
	PORT MAP (Z0 => UQVN_N90, A0 => UQVN_N86, A1 => UQVN_N85, A2 => UQVN_N84, 
	A3 => UQVN_N83, A4 => UQVN_N82, A5 => UQVN_N81, A6 => UQVN_N80, 
	A7 => UQVN_N79, A8 => UQVN_N78, A9 => UQVN_N77, A10 => UQVN_N76, 
	A11 => UQVN_N75);
UQVB_B112 : OR3
	PORT MAP (Z0 => UQVN_N88, A0 => UQVN_N87, A1 => UQVN_N89, A2 => UQVN_N90);
UQVB_B113 : INV
	PORT MAP (ZN0 => UQVN_N140, A0 => UQVN_N235);
UQVB_B114 : INV
	PORT MAP (ZN0 => UQVN_N138, A0 => B7);
UQVB_B115 : INV
	PORT MAP (ZN0 => UQVN_N139, A0 => B8);
UQVB_B116 : INV
	PORT MAP (ZN0 => UQVN_N134, A0 => A6);
UQVB_B117 : AND2
	PORT MAP (Z0 => UQVN_N98, A0 => UQVN_N137, A1 => UQVN_N235);
UQVB_B118 : AND2
	PORT MAP (Z0 => UQVN_N99, A0 => B6, A1 => UQVN_N140);
UQVB_B119 : OR2
	PORT MAP (Z0 => UQVN_N100, A0 => UQVN_N98, A1 => UQVN_N99);
UQVB_B120 : LXOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N100);
UQVB_B121 : AND3
	PORT MAP (Z0 => UQVN_N106, A0 => UQVN_N134, A1 => B7, A2 => UQVN_N137);
UQVB_B122 : AND3
	PORT MAP (Z0 => UQVN_N102, A0 => UQVN_N138, A1 => B6, A2 => UQVN_N235);
UQVB_B123 : AND3
	PORT MAP (Z0 => UQVN_N101, A0 => A6, A1 => UQVN_N138, A2 => UQVN_N235);
UQVB_B124 : AND3
	PORT MAP (Z0 => UQVN_N103, A0 => B7, A1 => UQVN_N137, A2 => UQVN_N140);
UQVB_B125 : AND3
	PORT MAP (Z0 => UQVN_N104, A0 => UQVN_N134, A1 => B7, A2 => UQVN_N140);
UQVB_B126 : OR6
	PORT MAP (Z0 => UQVN_N107, A0 => UQVN_N104, A1 => UQVN_N103, A2 => UQVN_N101, 
	A3 => UQVN_N102, A4 => UQVN_N106, A5 => UQVN_N105);
UQVB_B127 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N107);
UQVB_B128 : AND3
	PORT MAP (Z0 => UQVN_N105, A0 => A6, A1 => UQVN_N138, A2 => B6);
UQVB_B129 : AND4
	PORT MAP (Z0 => UQVN_N111, A0 => A6, A1 => A7, A2 => A8, 
	A3 => B6);
UQVB_B130 : AND3
	PORT MAP (Z0 => UQVN_N110, A0 => A7, A1 => A8, A2 => B7);
UQVB_B131 : AND4
	PORT MAP (Z0 => UQVN_N109, A0 => A6, A1 => A8, A2 => B6, 
	A3 => B7);
UQVB_B132 : AND2
	PORT MAP (Z0 => UQVN_N108, A0 => A8, A1 => B8);
UQVB_B133 : AND4
	PORT MAP (Z0 => UQVN_N112, A0 => A6, A1 => A7, A2 => B6, 
	A3 => B8);
UQVB_B134 : AND3
	PORT MAP (Z0 => UQVN_N113, A0 => A7, A1 => B7, A2 => B8);
UQVB_B135 : AND4
	PORT MAP (Z0 => UQVN_N114, A0 => A6, A1 => B6, A2 => B7, 
	A3 => B8);
UQVB_B136 : OR7
	PORT MAP (Z0 => G678, A0 => UQVN_N111, A1 => UQVN_N110, A2 => UQVN_N109, 
	A3 => UQVN_N108, A4 => UQVN_N112, A5 => UQVN_N113, A6 => UQVN_N114);
UQVB_B137 : AND2
	PORT MAP (Z0 => UQVN_N117, A0 => UQVN_N134, A1 => UQVN_N137);
UQVB_B138 : AND2
	PORT MAP (Z0 => UQVN_N115, A0 => UQVN_N135, A1 => UQVN_N138);
UQVB_B139 : AND2
	PORT MAP (Z0 => UQVN_N116, A0 => UQVN_N136, A1 => UQVN_N139);
UQVB_B140 : NOR3
	PORT MAP (ZN0 => P678, A0 => UQVN_N117, A1 => UQVN_N115, A2 => UQVN_N116);
UQVB_B141 : INV
	PORT MAP (ZN0 => UQVN_N137, A0 => B6);
UQVB_B142 : INV
	PORT MAP (ZN0 => UQVN_N135, A0 => A7);
UQVB_B143 : INV
	PORT MAP (ZN0 => UQVN_N136, A0 => A8);
UQVB_B144 : LXOR2
	PORT MAP (Z0 => Z8, A0 => A8, A1 => UQVN_N131);
UQVB_B145 : AND4
	PORT MAP (Z0 => UQVN_N130, A0 => UQVN_N137, A1 => UQVN_N138, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B146 : AND4
	PORT MAP (Z0 => UQVN_N132, A0 => UQVN_N134, A1 => UQVN_N138, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B147 : AND4
	PORT MAP (Z0 => UQVN_N129, A0 => UQVN_N135, A1 => UQVN_N137, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B148 : AND4
	PORT MAP (Z0 => UQVN_N128, A0 => UQVN_N134, A1 => UQVN_N135, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B149 : AND4
	PORT MAP (Z0 => UQVN_N127, A0 => B6, A1 => B7, A2 => UQVN_N139, 
	A3 => UQVN_N235);
UQVB_B150 : AND4
	PORT MAP (Z0 => UQVN_N126, A0 => A6, A1 => B7, A2 => UQVN_N139, 
	A3 => UQVN_N235);
UQVB_B151 : AND4
	PORT MAP (Z0 => UQVN_N125, A0 => A7, A1 => B6, A2 => UQVN_N139, 
	A3 => UQVN_N235);
UQVB_B152 : AND4
	PORT MAP (Z0 => UQVN_N124, A0 => A6, A1 => A7, A2 => UQVN_N139, 
	A3 => UQVN_N235);
UQVB_B153 : AND4
	PORT MAP (Z0 => UQVN_N123, A0 => A6, A1 => B6, A2 => B7, 
	A3 => UQVN_N139);
UQVB_B154 : AND3
	PORT MAP (Z0 => UQVN_N122, A0 => A7, A1 => B7, A2 => UQVN_N139);
UQVB_B155 : AND4
	PORT MAP (Z0 => UQVN_N121, A0 => A6, A1 => A7, A2 => B6, 
	A3 => UQVN_N139);
UQVB_B156 : AND4
	PORT MAP (Z0 => UQVN_N120, A0 => UQVN_N134, A1 => UQVN_N137, A2 => UQVN_N138, 
	A3 => B8);
UQVB_B157 : AND3
	PORT MAP (Z0 => UQVN_N119, A0 => UQVN_N135, A1 => UQVN_N138, A2 => B8);
UQVB_B158 : AND4
	PORT MAP (Z0 => UQVN_N118, A0 => UQVN_N134, A1 => UQVN_N135, A2 => UQVN_N137, 
	A3 => B8);
UQVB_B159 : OR12
	PORT MAP (Z0 => UQVN_N133, A0 => UQVN_N129, A1 => UQVN_N128, A2 => UQVN_N127, 
	A3 => UQVN_N126, A4 => UQVN_N125, A5 => UQVN_N124, A6 => UQVN_N123, 
	A7 => UQVN_N122, A8 => UQVN_N121, A9 => UQVN_N120, A10 => UQVN_N119, 
	A11 => UQVN_N118);
UQVB_B160 : OR3
	PORT MAP (Z0 => UQVN_N131, A0 => UQVN_N130, A1 => UQVN_N132, A2 => UQVN_N133);
UQVB_B161 : INV
	PORT MAP (ZN0 => UQVN_N183, A0 => UQVN_N236);
UQVB_B162 : INV
	PORT MAP (ZN0 => UQVN_N181, A0 => B10);
UQVB_B163 : INV
	PORT MAP (ZN0 => UQVN_N182, A0 => B11);
UQVB_B164 : INV
	PORT MAP (ZN0 => UQVN_N177, A0 => A9);
UQVB_B165 : AND2
	PORT MAP (Z0 => UQVN_N141, A0 => UQVN_N180, A1 => UQVN_N236);
UQVB_B166 : AND2
	PORT MAP (Z0 => UQVN_N142, A0 => B9, A1 => UQVN_N183);
UQVB_B167 : OR2
	PORT MAP (Z0 => UQVN_N143, A0 => UQVN_N141, A1 => UQVN_N142);
UQVB_B168 : LXOR2
	PORT MAP (Z0 => Z9, A0 => A9, A1 => UQVN_N143);
UQVB_B169 : AND3
	PORT MAP (Z0 => UQVN_N149, A0 => UQVN_N177, A1 => B10, A2 => UQVN_N180);
UQVB_B170 : AND3
	PORT MAP (Z0 => UQVN_N145, A0 => UQVN_N181, A1 => B9, A2 => UQVN_N236);
UQVB_B171 : AND3
	PORT MAP (Z0 => UQVN_N144, A0 => A9, A1 => UQVN_N181, A2 => UQVN_N236);
UQVB_B172 : AND3
	PORT MAP (Z0 => UQVN_N146, A0 => B10, A1 => UQVN_N180, A2 => UQVN_N183);
UQVB_B173 : AND3
	PORT MAP (Z0 => UQVN_N147, A0 => UQVN_N177, A1 => B10, A2 => UQVN_N183);
UQVB_B174 : OR6
	PORT MAP (Z0 => UQVN_N150, A0 => UQVN_N147, A1 => UQVN_N146, A2 => UQVN_N144, 
	A3 => UQVN_N145, A4 => UQVN_N149, A5 => UQVN_N148);
UQVB_B175 : LXOR2
	PORT MAP (Z0 => Z10, A0 => A10, A1 => UQVN_N150);
UQVB_B176 : AND3
	PORT MAP (Z0 => UQVN_N148, A0 => A9, A1 => UQVN_N181, A2 => B9);
UQVB_B177 : AND4
	PORT MAP (Z0 => UQVN_N154, A0 => A9, A1 => A10, A2 => A11, 
	A3 => B9);
UQVB_B178 : AND3
	PORT MAP (Z0 => UQVN_N153, A0 => A10, A1 => A11, A2 => B10);
UQVB_B179 : AND4
	PORT MAP (Z0 => UQVN_N152, A0 => A9, A1 => A11, A2 => B9, 
	A3 => B10);
UQVB_B180 : AND2
	PORT MAP (Z0 => UQVN_N151, A0 => A11, A1 => B11);
UQVB_B181 : AND4
	PORT MAP (Z0 => UQVN_N155, A0 => A9, A1 => A10, A2 => B9, 
	A3 => B11);
UQVB_B182 : AND3
	PORT MAP (Z0 => UQVN_N156, A0 => A10, A1 => B10, A2 => B11);
UQVB_B183 : AND4
	PORT MAP (Z0 => UQVN_N157, A0 => A9, A1 => B9, A2 => B10, 
	A3 => B11);
UQVB_B184 : OR7
	PORT MAP (Z0 => G911, A0 => UQVN_N154, A1 => UQVN_N153, A2 => UQVN_N152, 
	A3 => UQVN_N151, A4 => UQVN_N155, A5 => UQVN_N156, A6 => UQVN_N157);
UQVB_B185 : AND2
	PORT MAP (Z0 => UQVN_N160, A0 => UQVN_N177, A1 => UQVN_N180);
UQVB_B186 : AND2
	PORT MAP (Z0 => UQVN_N158, A0 => UQVN_N178, A1 => UQVN_N181);
UQVB_B187 : AND2
	PORT MAP (Z0 => UQVN_N159, A0 => UQVN_N179, A1 => UQVN_N182);
UQVB_B188 : NOR3
	PORT MAP (ZN0 => P911, A0 => UQVN_N160, A1 => UQVN_N158, A2 => UQVN_N159);
UQVB_B189 : INV
	PORT MAP (ZN0 => UQVN_N180, A0 => B9);
UQVB_B190 : INV
	PORT MAP (ZN0 => UQVN_N178, A0 => A10);
UQVB_B191 : INV
	PORT MAP (ZN0 => UQVN_N179, A0 => A11);
UQVB_B192 : LXOR2
	PORT MAP (Z0 => Z11, A0 => A11, A1 => UQVN_N174);
UQVB_B193 : AND4
	PORT MAP (Z0 => UQVN_N173, A0 => UQVN_N180, A1 => UQVN_N181, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B194 : AND4
	PORT MAP (Z0 => UQVN_N175, A0 => UQVN_N177, A1 => UQVN_N181, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B195 : AND4
	PORT MAP (Z0 => UQVN_N172, A0 => UQVN_N178, A1 => UQVN_N180, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B196 : AND4
	PORT MAP (Z0 => UQVN_N171, A0 => UQVN_N177, A1 => UQVN_N178, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B197 : AND4
	PORT MAP (Z0 => UQVN_N170, A0 => B9, A1 => B10, A2 => UQVN_N182, 
	A3 => UQVN_N236);
UQVB_B198 : AND4
	PORT MAP (Z0 => UQVN_N169, A0 => A9, A1 => B10, A2 => UQVN_N182, 
	A3 => UQVN_N236);
UQVB_B199 : AND4
	PORT MAP (Z0 => UQVN_N168, A0 => A10, A1 => B9, A2 => UQVN_N182, 
	A3 => UQVN_N236);
UQVB_B200 : AND4
	PORT MAP (Z0 => UQVN_N167, A0 => A9, A1 => A10, A2 => UQVN_N182, 
	A3 => UQVN_N236);
UQVB_B201 : AND4
	PORT MAP (Z0 => UQVN_N166, A0 => A9, A1 => B9, A2 => B10, 
	A3 => UQVN_N182);
UQVB_B202 : AND3
	PORT MAP (Z0 => UQVN_N165, A0 => A10, A1 => B10, A2 => UQVN_N182);
UQVB_B203 : AND4
	PORT MAP (Z0 => UQVN_N164, A0 => A9, A1 => A10, A2 => B9, 
	A3 => UQVN_N182);
UQVB_B204 : AND4
	PORT MAP (Z0 => UQVN_N163, A0 => UQVN_N177, A1 => UQVN_N180, A2 => UQVN_N181, 
	A3 => B11);
UQVB_B205 : AND3
	PORT MAP (Z0 => UQVN_N162, A0 => UQVN_N178, A1 => UQVN_N181, A2 => B11);
UQVB_B206 : AND4
	PORT MAP (Z0 => UQVN_N161, A0 => UQVN_N177, A1 => UQVN_N178, A2 => UQVN_N180, 
	A3 => B11);
UQVB_B207 : OR12
	PORT MAP (Z0 => UQVN_N176, A0 => UQVN_N172, A1 => UQVN_N171, A2 => UQVN_N170, 
	A3 => UQVN_N169, A4 => UQVN_N168, A5 => UQVN_N167, A6 => UQVN_N166, 
	A7 => UQVN_N165, A8 => UQVN_N164, A9 => UQVN_N163, A10 => UQVN_N162, 
	A11 => UQVN_N161);
UQVB_B208 : OR3
	PORT MAP (Z0 => UQVN_N174, A0 => UQVN_N173, A1 => UQVN_N175, A2 => UQVN_N176);
UQVB_B209 : INV
	PORT MAP (ZN0 => UQVN_N226, A0 => UQVN_N237);
UQVB_B210 : INV
	PORT MAP (ZN0 => UQVN_N224, A0 => B13);
UQVB_B211 : INV
	PORT MAP (ZN0 => UQVN_N225, A0 => B14);
UQVB_B212 : INV
	PORT MAP (ZN0 => UQVN_N220, A0 => A12);
UQVB_B213 : AND2
	PORT MAP (Z0 => UQVN_N184, A0 => UQVN_N223, A1 => UQVN_N237);
UQVB_B214 : AND2
	PORT MAP (Z0 => UQVN_N185, A0 => B12, A1 => UQVN_N226);
UQVB_B215 : OR2
	PORT MAP (Z0 => UQVN_N186, A0 => UQVN_N184, A1 => UQVN_N185);
UQVB_B216 : LXOR2
	PORT MAP (Z0 => Z12, A0 => A12, A1 => UQVN_N186);
UQVB_B217 : AND3
	PORT MAP (Z0 => UQVN_N192, A0 => UQVN_N220, A1 => B13, A2 => UQVN_N223);
UQVB_B218 : AND3
	PORT MAP (Z0 => UQVN_N188, A0 => UQVN_N224, A1 => B12, A2 => UQVN_N237);
UQVB_B219 : AND3
	PORT MAP (Z0 => UQVN_N187, A0 => A12, A1 => UQVN_N224, A2 => UQVN_N237);
UQVB_B220 : AND3
	PORT MAP (Z0 => UQVN_N189, A0 => B13, A1 => UQVN_N223, A2 => UQVN_N226);
UQVB_B221 : AND3
	PORT MAP (Z0 => UQVN_N190, A0 => UQVN_N220, A1 => B13, A2 => UQVN_N226);
UQVB_B222 : OR6
	PORT MAP (Z0 => UQVN_N193, A0 => UQVN_N190, A1 => UQVN_N189, A2 => UQVN_N187, 
	A3 => UQVN_N188, A4 => UQVN_N192, A5 => UQVN_N191);
UQVB_B223 : LXOR2
	PORT MAP (Z0 => Z13, A0 => A13, A1 => UQVN_N193);
UQVB_B224 : AND3
	PORT MAP (Z0 => UQVN_N191, A0 => A12, A1 => UQVN_N224, A2 => B12);
UQVB_B225 : AND4
	PORT MAP (Z0 => UQVN_N197, A0 => A12, A1 => A13, A2 => A14, 
	A3 => B12);
UQVB_B226 : AND3
	PORT MAP (Z0 => UQVN_N196, A0 => A13, A1 => A14, A2 => B13);
UQVB_B227 : AND4
	PORT MAP (Z0 => UQVN_N195, A0 => A12, A1 => A14, A2 => B12, 
	A3 => B13);
UQVB_B228 : AND2
	PORT MAP (Z0 => UQVN_N194, A0 => A14, A1 => B14);
UQVB_B229 : AND4
	PORT MAP (Z0 => UQVN_N198, A0 => A12, A1 => A13, A2 => B12, 
	A3 => B14);
UQVB_B230 : AND3
	PORT MAP (Z0 => UQVN_N199, A0 => A13, A1 => B13, A2 => B14);
UQVB_B231 : AND4
	PORT MAP (Z0 => UQVN_N200, A0 => A12, A1 => B12, A2 => B13, 
	A3 => B14);
UQVB_B232 : OR7
	PORT MAP (Z0 => G1214, A0 => UQVN_N197, A1 => UQVN_N196, A2 => UQVN_N195, 
	A3 => UQVN_N194, A4 => UQVN_N198, A5 => UQVN_N199, A6 => UQVN_N200);
UQVB_B233 : AND2
	PORT MAP (Z0 => UQVN_N203, A0 => UQVN_N220, A1 => UQVN_N223);
UQVB_B234 : AND2
	PORT MAP (Z0 => UQVN_N201, A0 => UQVN_N221, A1 => UQVN_N224);
UQVB_B235 : AND2
	PORT MAP (Z0 => UQVN_N202, A0 => UQVN_N222, A1 => UQVN_N225);
UQVB_B236 : NOR3
	PORT MAP (ZN0 => P1214, A0 => UQVN_N203, A1 => UQVN_N201, A2 => UQVN_N202);
UQVB_B237 : INV
	PORT MAP (ZN0 => UQVN_N223, A0 => B12);
UQVB_B238 : INV
	PORT MAP (ZN0 => UQVN_N221, A0 => A13);
UQVB_B239 : INV
	PORT MAP (ZN0 => UQVN_N222, A0 => A14);
UQVB_B240 : LXOR2
	PORT MAP (Z0 => Z14, A0 => A14, A1 => UQVN_N217);
UQVB_B241 : AND4
	PORT MAP (Z0 => UQVN_N216, A0 => UQVN_N223, A1 => UQVN_N224, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B242 : AND4
	PORT MAP (Z0 => UQVN_N218, A0 => UQVN_N220, A1 => UQVN_N224, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B243 : AND4
	PORT MAP (Z0 => UQVN_N215, A0 => UQVN_N221, A1 => UQVN_N223, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B244 : AND4
	PORT MAP (Z0 => UQVN_N214, A0 => UQVN_N220, A1 => UQVN_N221, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B245 : AND4
	PORT MAP (Z0 => UQVN_N213, A0 => B12, A1 => B13, A2 => UQVN_N225, 
	A3 => UQVN_N237);
UQVB_B246 : AND4
	PORT MAP (Z0 => UQVN_N212, A0 => A12, A1 => B13, A2 => UQVN_N225, 
	A3 => UQVN_N237);
UQVB_B247 : AND4
	PORT MAP (Z0 => UQVN_N211, A0 => A13, A1 => B12, A2 => UQVN_N225, 
	A3 => UQVN_N237);
UQVB_B248 : AND4
	PORT MAP (Z0 => UQVN_N210, A0 => A12, A1 => A13, A2 => UQVN_N225, 
	A3 => UQVN_N237);
UQVB_B249 : AND4
	PORT MAP (Z0 => UQVN_N209, A0 => A12, A1 => B12, A2 => B13, 
	A3 => UQVN_N225);
UQVB_B250 : AND3
	PORT MAP (Z0 => UQVN_N208, A0 => A13, A1 => B13, A2 => UQVN_N225);
UQVB_B251 : AND4
	PORT MAP (Z0 => UQVN_N207, A0 => A12, A1 => A13, A2 => B12, 
	A3 => UQVN_N225);
UQVB_B252 : AND4
	PORT MAP (Z0 => UQVN_N206, A0 => UQVN_N220, A1 => UQVN_N223, A2 => UQVN_N224, 
	A3 => B14);
UQVB_B253 : AND3
	PORT MAP (Z0 => UQVN_N205, A0 => UQVN_N221, A1 => UQVN_N224, A2 => B14);
UQVB_B254 : AND4
	PORT MAP (Z0 => UQVN_N204, A0 => UQVN_N220, A1 => UQVN_N221, A2 => UQVN_N223, 
	A3 => B14);
UQVB_B255 : OR12
	PORT MAP (Z0 => UQVN_N219, A0 => UQVN_N215, A1 => UQVN_N214, A2 => UQVN_N213, 
	A3 => UQVN_N212, A4 => UQVN_N211, A5 => UQVN_N210, A6 => UQVN_N209, 
	A7 => UQVN_N208, A8 => UQVN_N207, A9 => UQVN_N206, A10 => UQVN_N205, 
	A11 => UQVN_N204);
UQVB_B256 : OR3
	PORT MAP (Z0 => UQVN_N217, A0 => UQVN_N216, A1 => UQVN_N218, A2 => UQVN_N219);
UQVB_B257 : AND2
	PORT MAP (Z0 => UQVN_N228, A0 => UQVN_N234, A1 => UQVN_N238);
UQVB_B258 : AND2
	PORT MAP (Z0 => UQVN_N229, A0 => B15, A1 => UQVN_N227);
UQVB_B259 : OR2
	PORT MAP (Z0 => UQVN_N230, A0 => UQVN_N229, A1 => UQVN_N228);
UQVB_B260 : XOR2
	PORT MAP (Z0 => Z15, A0 => A15, A1 => UQVN_N230);
UQVB_B261 : INV
	PORT MAP (ZN0 => UQVN_N234, A0 => B15);
UQVB_B262 : INV
	PORT MAP (ZN0 => UQVN_N227, A0 => UQVN_N238);
UQVB_B263 : AND2
	PORT MAP (Z0 => UQVN_N231, A0 => UQVN_N238, A1 => B15);
UQVB_B264 : AND2
	PORT MAP (Z0 => UQVN_N232, A0 => UQVN_N238, A1 => A15);
UQVB_B265 : AND2
	PORT MAP (Z0 => UQVN_N233, A0 => B15, A1 => A15);
UQVB_B266 : OR3
	PORT MAP (Z0 => CO, A0 => UQVN_N231, A1 => UQVN_N232, A2 => UQVN_N233);
END lattice_arch;
-- VHDL netlist for ADDF2
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDF2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDF2;


ARCHITECTURE lattice_arch OF ADDF2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => CI);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => CI, A1 => A1, A2 => A0);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => CI, A1 => A1, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => CI, A1 => A0, A2 => B1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => CI, A1 => B1, A2 => B0);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A1, A1 => A0, A2 => B0);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A0, A1 => B1, A2 => B0);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => A1, A1 => B1);
UQVB_B9 : OR7
	PORT MAP (Z0 => CO, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N5, A5 => UQVN_N7, A6 => UQVN_N6);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N18, A1 => B1, A2 => UQVN_N21);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B1, A1 => UQVN_N19, A2 => UQVN_N21);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => A0, A1 => UQVN_N20, A2 => CI);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N20, A1 => B0, A2 => CI);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N18, A1 => B1, A2 => UQVN_N19);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A0, A1 => UQVN_N20, A2 => B0);
UQVB_B16 : OR6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N12, A5 => UQVN_N13);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N14);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => B0);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => B1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => A0);
UQVB_B21 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N15);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => CI, A1 => UQVN_N19);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N16, A1 => UQVN_N17);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N21, A1 => B0);
END lattice_arch;
-- VHDL netlist for ADDF4
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDF4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDF4;


ARCHITECTURE lattice_arch OF ADDF4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => CI);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => CI, A1 => A1, A2 => A0);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => CI, A1 => A1, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => CI, A1 => A0, A2 => B1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => CI, A1 => B1, A2 => B0);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A1, A1 => A0, A2 => B0);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A0, A1 => B1, A2 => B0);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => A1, A1 => B1);
UQVB_B9 : OR7
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N5, A5 => UQVN_N7, A6 => UQVN_N6);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N18, A1 => B1, A2 => UQVN_N21);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B1, A1 => UQVN_N19, A2 => UQVN_N21);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => A0, A1 => UQVN_N20, A2 => CI);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N20, A1 => B0, A2 => CI);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N18, A1 => B1, A2 => UQVN_N19);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A0, A1 => UQVN_N20, A2 => B0);
UQVB_B16 : OR6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N12, A5 => UQVN_N13);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N14);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => B0);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => B1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => A0);
UQVB_B21 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N15);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => CI, A1 => UQVN_N19);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N16, A1 => UQVN_N17);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N21, A1 => B0);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => UQVN_N43);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N43, A1 => A3, A2 => A2);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N43, A1 => A3, A2 => B2);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N43, A1 => A2, A2 => B3);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N43, A1 => B3, A2 => B2);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => A3, A1 => A2, A2 => B2);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => A2, A1 => B3, A2 => B2);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => A3, A1 => B3);
UQVB_B33 : OR7
	PORT MAP (Z0 => CO, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N22, 
	A3 => UQVN_N25, A4 => UQVN_N26, A5 => UQVN_N28, A6 => UQVN_N27);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N39, A1 => B3, A2 => UQVN_N42);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => B3, A1 => UQVN_N40, A2 => UQVN_N42);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => A2, A1 => UQVN_N41, A2 => UQVN_N43);
UQVB_B37 : AND3
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N41, A1 => B2, A2 => UQVN_N43);
UQVB_B38 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N39, A1 => B3, A2 => UQVN_N40);
UQVB_B39 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => A2, A1 => UQVN_N41, A2 => B2);
UQVB_B40 : OR6
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N29, A1 => UQVN_N30, A2 => UQVN_N31, 
	A3 => UQVN_N32, A4 => UQVN_N33, A5 => UQVN_N34);
UQVB_B41 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N35);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => B2);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B3);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A2);
UQVB_B45 : XOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N36);
UQVB_B46 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N43, A1 => UQVN_N40);
UQVB_B47 : OR2
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N37, A1 => UQVN_N38);
UQVB_B48 : AND2
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N42, A1 => B2);
END lattice_arch;
-- VHDL netlist for ADDF8
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDF8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDF8;


ARCHITECTURE lattice_arch OF ADDF8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, G0, G1, G2,
	 G3, G4, G5, G6,
	 G7, P0, P1, P2,
	 P3, P4, P5, P6,
	 P7 : std_logic;


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : XOR2
	PORT MAP (Z0 => P7, A0 => A7, A1 => B7);
UQVB_B2 : XOR2
	PORT MAP (Z0 => P6, A0 => A6, A1 => B6);
UQVB_B3 : XOR2
	PORT MAP (Z0 => P5, A0 => A5, A1 => B5);
UQVB_B4 : XOR2
	PORT MAP (Z0 => P4, A0 => A4, A1 => B4);
UQVB_B5 : XOR2
	PORT MAP (Z0 => P3, A0 => A3, A1 => B3);
UQVB_B6 : XOR2
	PORT MAP (Z0 => P2, A0 => A2, A1 => B2);
UQVB_B7 : XOR2
	PORT MAP (Z0 => P1, A0 => A1, A1 => B1);
UQVB_B8 : XOR2
	PORT MAP (Z0 => P0, A0 => A0, A1 => B0);
UQVB_B9 : AND2
	PORT MAP (Z0 => G7, A0 => A7, A1 => B7);
UQVB_B10 : AND2
	PORT MAP (Z0 => G6, A0 => A6, A1 => B6);
UQVB_B11 : AND2
	PORT MAP (Z0 => G5, A0 => A5, A1 => B5);
UQVB_B12 : AND2
	PORT MAP (Z0 => G4, A0 => A4, A1 => B4);
UQVB_B13 : AND2
	PORT MAP (Z0 => G3, A0 => A3, A1 => B3);
UQVB_B14 : AND2
	PORT MAP (Z0 => G2, A0 => A2, A1 => B2);
UQVB_B15 : AND2
	PORT MAP (Z0 => G1, A0 => A1, A1 => B1);
UQVB_B16 : AND2
	PORT MAP (Z0 => G0, A0 => A0, A1 => B0);
UQVB_B17 : AND8
	PORT MAP (Z0 => UQVN_N11, A0 => G0, A1 => P1, A2 => P2, 
	A3 => P3, A4 => P4, A5 => P5, A6 => P6, 
	A7 => P7);
UQVB_B18 : OR6
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N5, A5 => G4);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N6, A1 => P5);
UQVB_B20 : AND7
	PORT MAP (Z0 => UQVN_N10, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4, A4 => P5, A5 => P6, A6 => P7);
UQVB_B21 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N15, A1 => UQVN_N14, A2 => UQVN_N17, 
	A3 => UQVN_N16, A4 => G7);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => G0, A1 => P1);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => CI, A1 => P0, A2 => P1);
UQVB_B24 : OR3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N7, A1 => UQVN_N8, A2 => G1);
UQVB_B25 : AND9
	PORT MAP (Z0 => UQVN_N13, A0 => CI, A1 => P0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4, A6 => P5, 
	A7 => P6, A8 => P7);
UQVB_B26 : LXOR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N9, A1 => P2);
UQVB_B27 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => G2, A1 => P3, A2 => P4, 
	A3 => P5, A4 => P6, A5 => P7);
UQVB_B28 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => G3, A1 => P4, A2 => P5, 
	A3 => P6, A4 => P7);
UQVB_B29 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => G6, A1 => P7);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => G5, A1 => P6, A2 => P7);
UQVB_B31 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => G4, A1 => P5, A2 => P6, 
	A3 => P7);
UQVB_B32 : OR4
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N13, A1 => UQVN_N11, A2 => UQVN_N10, 
	A3 => UQVN_N12);
UQVB_B33 : OR2
	PORT MAP (Z0 => CO, A0 => UQVN_N19, A1 => UQVN_N18);
UQVB_B34 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => CI, A1 => P0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => G0, A1 => P1, A2 => P2, 
	A3 => P3, A4 => P4);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4);
UQVB_B37 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => G2, A1 => P3, A2 => P4);
UQVB_B38 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => G3, A1 => P4);
UQVB_B39 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => CI, A1 => P0);
UQVB_B40 : OR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N31, A1 => G0);
UQVB_B41 : OR2
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N21, A1 => UQVN_N20);
UQVB_B42 : LXOR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N30, A1 => P1);
UQVB_B43 : XOR2
	PORT MAP (Z0 => Z0, A0 => CI, A1 => P0);
UQVB_B44 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => G5, A1 => P6);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => G4, A1 => P5, A2 => P6);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => G3, A1 => P4, A2 => P5, 
	A3 => P6);
UQVB_B47 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => G2, A1 => P3, A2 => P4, 
	A3 => P5, A4 => P6);
UQVB_B48 : AND6
	PORT MAP (Z0 => UQVN_N22, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4, A4 => P5, A5 => P6);
UQVB_B49 : AND7
	PORT MAP (Z0 => UQVN_N23, A0 => G0, A1 => P1, A2 => P2, 
	A3 => P3, A4 => P4, A5 => P5, A6 => P6);
UQVB_B50 : AND8
	PORT MAP (Z0 => UQVN_N25, A0 => CI, A1 => P0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4, A6 => P5, 
	A7 => P6);
UQVB_B51 : OR5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N25, A1 => UQVN_N23, A2 => UQVN_N22, 
	A3 => UQVN_N24, A4 => UQVN_N27);
UQVB_B52 : OR3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N26, A1 => UQVN_N28, A2 => G6);
UQVB_B53 : LXOR2
	PORT MAP (Z0 => Z7, A0 => UQVN_N29, A1 => P7);
UQVB_B54 : AND2
	PORT MAP (Z0 => UQVN_N46, A0 => G2, A1 => P3);
UQVB_B55 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => G1, A1 => P2, A2 => P3);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N47, A0 => G0, A1 => P1, A2 => P2, 
	A3 => P3);
UQVB_B57 : AND5
	PORT MAP (Z0 => UQVN_N48, A0 => CI, A1 => P0, A2 => P1, 
	A3 => P2, A4 => P3);
UQVB_B58 : OR5
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N48, A1 => UQVN_N47, A2 => UQVN_N45, 
	A3 => UQVN_N46, A4 => G3);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N32, A1 => P3);
UQVB_B60 : AND2
	PORT MAP (Z0 => UQVN_N35, A0 => G1, A1 => P2);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => G0, A1 => P1, A2 => P2);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => CI, A1 => P0, A2 => P1, 
	A3 => P2);
UQVB_B63 : OR4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N33, A1 => UQVN_N34, A2 => UQVN_N35, 
	A3 => G2);
UQVB_B64 : OR2
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N37, A1 => UQVN_N36);
UQVB_B65 : OR4
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N41, A1 => UQVN_N39, A2 => UQVN_N38, 
	A3 => UQVN_N40);
UQVB_B66 : LXOR2
	PORT MAP (Z0 => Z4, A0 => UQVN_N44, A1 => P4);
UQVB_B67 : AND2
	PORT MAP (Z0 => UQVN_N42, A0 => G4, A1 => P5);
UQVB_B68 : AND3
	PORT MAP (Z0 => UQVN_N43, A0 => G3, A1 => P4, A2 => P5);
UQVB_B69 : AND4
	PORT MAP (Z0 => UQVN_N40, A0 => G2, A1 => P3, A2 => P4, 
	A3 => P5);
UQVB_B70 : AND5
	PORT MAP (Z0 => UQVN_N38, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4, A4 => P5);
UQVB_B71 : AND6
	PORT MAP (Z0 => UQVN_N39, A0 => G0, A1 => P1, A2 => P2, 
	A3 => P3, A4 => P4, A5 => P5);
UQVB_B72 : AND7
	PORT MAP (Z0 => UQVN_N41, A0 => CI, A1 => P0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4, A6 => P5);
UQVB_B73 : OR3
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N43, A1 => UQVN_N42, A2 => G5);
UQVB_B74 : LXOR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N49, A1 => P6);
END lattice_arch;
-- VHDL netlist for ADDF8A
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDF8A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDF8A;


ARCHITECTURE lattice_arch OF ADDF8A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 G012, G345, P012, P345 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => CI);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B2);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => A0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N40, A1 => CI);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => UQVN_N43);
UQVB_B7 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N3);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N37, A1 => B1, A2 => UQVN_N40);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N41, A1 => B0, A2 => CI);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => A0, A1 => UQVN_N41, A2 => CI);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B1, A1 => UQVN_N40, A2 => UQVN_N43);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N37, A1 => B1, A2 => UQVN_N43);
UQVB_B14 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N8);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => UQVN_N41, A2 => B0);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => A0, A1 => A1, A2 => A2, 
	A3 => B0);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A1, A1 => A2, A2 => B1);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => A0, A1 => A2, A2 => B0, 
	A3 => B1);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A2, A1 => B2);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B2);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => A1, A1 => B1, A2 => B2);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => A0, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B24 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16, A6 => UQVN_N17);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N37, A1 => UQVN_N40);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N38, A1 => UQVN_N41);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N39, A1 => UQVN_N42);
UQVB_B28 : NOR3
	PORT MAP (ZN0 => P012, A0 => UQVN_N20, A1 => UQVN_N18, A2 => UQVN_N19);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => B0);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A1);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A2);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N34);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N41, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N38, A1 => UQVN_N40, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N37, A1 => UQVN_N38, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => B0, A1 => B1, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => A0, A1 => B1, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A1, A1 => B0, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => A0, A1 => A1, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => A0, A1 => B0, A2 => B1, 
	A3 => UQVN_N42);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => A1, A1 => B1, A2 => UQVN_N42);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => A0, A1 => A1, A2 => B0, 
	A3 => UQVN_N42);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N37, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => B2);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N38, A1 => UQVN_N41, A2 => B2);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N37, A1 => UQVN_N38, A2 => UQVN_N40, 
	A3 => B2);
UQVB_B47 : OR12
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N28, A5 => UQVN_N27, A6 => UQVN_N26, 
	A7 => UQVN_N25, A8 => UQVN_N24, A9 => UQVN_N23, A10 => UQVN_N22, 
	A11 => UQVN_N21);
UQVB_B48 : OR3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N33, A1 => UQVN_N35, A2 => UQVN_N36);
UQVB_B49 : AND2
	PORT MAP (Z0 => UQVN_N44, A0 => P012, A1 => CI);
UQVB_B50 : OR2
	PORT MAP (Z0 => UQVN_N111, A0 => G012, A1 => UQVN_N44);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N87, A0 => UQVN_N111);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N85, A0 => B4);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N86, A0 => B5);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N81, A0 => A3);
UQVB_B55 : AND2
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N84, A1 => UQVN_N111);
UQVB_B56 : AND2
	PORT MAP (Z0 => UQVN_N46, A0 => B3, A1 => UQVN_N87);
UQVB_B57 : OR2
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N45, A1 => UQVN_N46);
UQVB_B58 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N47);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N81, A1 => B4, A2 => UQVN_N84);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N85, A1 => B3, A2 => UQVN_N111);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N48, A0 => A3, A1 => UQVN_N85, A2 => UQVN_N111);
UQVB_B62 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => B4, A1 => UQVN_N84, A2 => UQVN_N87);
UQVB_B63 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N81, A1 => B4, A2 => UQVN_N87);
UQVB_B64 : OR6
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N51, A1 => UQVN_N50, A2 => UQVN_N48, 
	A3 => UQVN_N49, A4 => UQVN_N53, A5 => UQVN_N52);
UQVB_B65 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N54);
UQVB_B66 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => A3, A1 => UQVN_N85, A2 => B3);
UQVB_B67 : AND4
	PORT MAP (Z0 => UQVN_N58, A0 => A3, A1 => A4, A2 => A5, 
	A3 => B3);
UQVB_B68 : AND3
	PORT MAP (Z0 => UQVN_N57, A0 => A4, A1 => A5, A2 => B4);
UQVB_B69 : AND4
	PORT MAP (Z0 => UQVN_N56, A0 => A3, A1 => A5, A2 => B3, 
	A3 => B4);
UQVB_B70 : AND2
	PORT MAP (Z0 => UQVN_N55, A0 => A5, A1 => B5);
UQVB_B71 : AND4
	PORT MAP (Z0 => UQVN_N59, A0 => A3, A1 => A4, A2 => B3, 
	A3 => B5);
UQVB_B72 : AND3
	PORT MAP (Z0 => UQVN_N60, A0 => A4, A1 => B4, A2 => B5);
UQVB_B73 : AND4
	PORT MAP (Z0 => UQVN_N61, A0 => A3, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B74 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N58, A1 => UQVN_N57, A2 => UQVN_N56, 
	A3 => UQVN_N55, A4 => UQVN_N59, A5 => UQVN_N60, A6 => UQVN_N61);
UQVB_B75 : AND2
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N81, A1 => UQVN_N84);
UQVB_B76 : AND2
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N82, A1 => UQVN_N85);
UQVB_B77 : AND2
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N83, A1 => UQVN_N86);
UQVB_B78 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N64, A1 => UQVN_N62, A2 => UQVN_N63);
UQVB_B79 : INV
	PORT MAP (ZN0 => UQVN_N84, A0 => B3);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N82, A0 => A4);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N83, A0 => A5);
UQVB_B82 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N78);
UQVB_B83 : AND4
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N84, A1 => UQVN_N85, A2 => B5, 
	A3 => UQVN_N87);
UQVB_B84 : AND4
	PORT MAP (Z0 => UQVN_N79, A0 => UQVN_N81, A1 => UQVN_N85, A2 => B5, 
	A3 => UQVN_N87);
UQVB_B85 : AND4
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N82, A1 => UQVN_N84, A2 => B5, 
	A3 => UQVN_N87);
UQVB_B86 : AND4
	PORT MAP (Z0 => UQVN_N75, A0 => UQVN_N81, A1 => UQVN_N82, A2 => B5, 
	A3 => UQVN_N87);
UQVB_B87 : AND4
	PORT MAP (Z0 => UQVN_N74, A0 => B3, A1 => B4, A2 => UQVN_N86, 
	A3 => UQVN_N111);
UQVB_B88 : AND4
	PORT MAP (Z0 => UQVN_N73, A0 => A3, A1 => B4, A2 => UQVN_N86, 
	A3 => UQVN_N111);
UQVB_B89 : AND4
	PORT MAP (Z0 => UQVN_N72, A0 => A4, A1 => B3, A2 => UQVN_N86, 
	A3 => UQVN_N111);
UQVB_B90 : AND4
	PORT MAP (Z0 => UQVN_N71, A0 => A3, A1 => A4, A2 => UQVN_N86, 
	A3 => UQVN_N111);
UQVB_B91 : AND4
	PORT MAP (Z0 => UQVN_N70, A0 => A3, A1 => B3, A2 => B4, 
	A3 => UQVN_N86);
UQVB_B92 : AND3
	PORT MAP (Z0 => UQVN_N69, A0 => A4, A1 => B4, A2 => UQVN_N86);
UQVB_B93 : AND4
	PORT MAP (Z0 => UQVN_N68, A0 => A3, A1 => A4, A2 => B3, 
	A3 => UQVN_N86);
UQVB_B94 : AND4
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N81, A1 => UQVN_N84, A2 => UQVN_N85, 
	A3 => B5);
UQVB_B95 : AND3
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N82, A1 => UQVN_N85, A2 => B5);
UQVB_B96 : AND4
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N81, A1 => UQVN_N82, A2 => UQVN_N84, 
	A3 => B5);
UQVB_B97 : OR12
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N76, A1 => UQVN_N75, A2 => UQVN_N74, 
	A3 => UQVN_N73, A4 => UQVN_N72, A5 => UQVN_N71, A6 => UQVN_N70, 
	A7 => UQVN_N69, A8 => UQVN_N68, A9 => UQVN_N67, A10 => UQVN_N66, 
	A11 => UQVN_N65);
UQVB_B98 : OR3
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N77, A1 => UQVN_N79, A2 => UQVN_N80);
UQVB_B99 : OR3
	PORT MAP (Z0 => UQVN_N112, A0 => G345, A1 => UQVN_N88, A2 => UQVN_N89);
UQVB_B100 : AND3
	PORT MAP (Z0 => UQVN_N89, A0 => P345, A1 => P012, A2 => CI);
UQVB_B101 : AND2
	PORT MAP (Z0 => UQVN_N88, A0 => P345, A1 => G012);
UQVB_B102 : INV
	PORT MAP (ZN0 => UQVN_N110, A0 => UQVN_N112);
UQVB_B103 : AND3
	PORT MAP (Z0 => UQVN_N92, A0 => UQVN_N112, A1 => A7, A2 => A6);
UQVB_B104 : AND3
	PORT MAP (Z0 => UQVN_N91, A0 => UQVN_N112, A1 => A7, A2 => B6);
UQVB_B105 : AND3
	PORT MAP (Z0 => UQVN_N90, A0 => UQVN_N112, A1 => A6, A2 => B7);
UQVB_B106 : AND3
	PORT MAP (Z0 => UQVN_N93, A0 => UQVN_N112, A1 => B7, A2 => B6);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N94, A0 => A7, A1 => A6, A2 => B6);
UQVB_B108 : AND3
	PORT MAP (Z0 => UQVN_N96, A0 => A6, A1 => B7, A2 => B6);
UQVB_B109 : AND2
	PORT MAP (Z0 => UQVN_N95, A0 => A7, A1 => B7);
UQVB_B110 : OR7
	PORT MAP (Z0 => CO, A0 => UQVN_N92, A1 => UQVN_N91, A2 => UQVN_N90, 
	A3 => UQVN_N93, A4 => UQVN_N94, A5 => UQVN_N96, A6 => UQVN_N95);
UQVB_B111 : AND3
	PORT MAP (Z0 => UQVN_N97, A0 => UQVN_N107, A1 => B7, A2 => UQVN_N110);
UQVB_B112 : AND3
	PORT MAP (Z0 => UQVN_N98, A0 => B7, A1 => UQVN_N108, A2 => UQVN_N110);
UQVB_B113 : AND3
	PORT MAP (Z0 => UQVN_N99, A0 => A6, A1 => UQVN_N109, A2 => UQVN_N112);
UQVB_B114 : AND3
	PORT MAP (Z0 => UQVN_N100, A0 => UQVN_N109, A1 => B6, A2 => UQVN_N112);
UQVB_B115 : AND3
	PORT MAP (Z0 => UQVN_N101, A0 => UQVN_N107, A1 => B7, A2 => UQVN_N108);
UQVB_B116 : AND3
	PORT MAP (Z0 => UQVN_N102, A0 => A6, A1 => UQVN_N109, A2 => B6);
UQVB_B117 : OR6
	PORT MAP (Z0 => UQVN_N103, A0 => UQVN_N97, A1 => UQVN_N98, A2 => UQVN_N99, 
	A3 => UQVN_N100, A4 => UQVN_N101, A5 => UQVN_N102);
UQVB_B118 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N103);
UQVB_B119 : INV
	PORT MAP (ZN0 => UQVN_N108, A0 => B6);
UQVB_B120 : INV
	PORT MAP (ZN0 => UQVN_N109, A0 => B7);
UQVB_B121 : INV
	PORT MAP (ZN0 => UQVN_N107, A0 => A6);
UQVB_B122 : XOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N104);
UQVB_B123 : AND2
	PORT MAP (Z0 => UQVN_N105, A0 => UQVN_N112, A1 => UQVN_N108);
UQVB_B124 : OR2
	PORT MAP (Z0 => UQVN_N104, A0 => UQVN_N105, A1 => UQVN_N106);
UQVB_B125 : AND2
	PORT MAP (Z0 => UQVN_N106, A0 => UQVN_N110, A1 => B6);
END lattice_arch;
-- VHDL netlist for ADDH1
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH1 IS 
    PORT (
        A0 : IN std_logic;
        B0 : IN std_logic;
        Z0 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDH1;


ARCHITECTURE lattice_arch OF ADDH1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N4, A1 => B0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N3, A1 => A0);
UQVB_B3 : AND2
	PORT MAP (Z0 => CO, A0 => B0, A1 => A0);
UQVB_B4 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => B0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
END lattice_arch;
-- VHDL netlist for ADDH16A
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH16A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B10 : IN std_logic;
        B11 : IN std_logic;
        B12 : IN std_logic;
        B13 : IN std_logic;
        B14 : IN std_logic;
        B15 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        B8 : IN std_logic;
        B9 : IN std_logic;
        CO : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z10 : OUT std_logic;
        Z11 : OUT std_logic;
        Z12 : OUT std_logic;
        Z13 : OUT std_logic;
        Z14 : OUT std_logic;
        Z15 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        Z8 : OUT std_logic;
        Z9 : OUT std_logic
    );
END ADDH16A;


ARCHITECTURE lattice_arch OF ADDH16A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 UQVN_N113, UQVN_N114, UQVN_N115, UQVN_N116,
	 UQVN_N117, UQVN_N118, UQVN_N119, UQVN_N120,
	 UQVN_N121, UQVN_N122, UQVN_N123, UQVN_N124,
	 UQVN_N125, UQVN_N126, UQVN_N127, UQVN_N128,
	 UQVN_N129, UQVN_N130, UQVN_N131, UQVN_N132,
	 UQVN_N133, UQVN_N134, UQVN_N135, UQVN_N136,
	 UQVN_N137, UQVN_N138, UQVN_N139, UQVN_N140,
	 UQVN_N141, UQVN_N142, UQVN_N143, UQVN_N144,
	 UQVN_N145, UQVN_N146, UQVN_N147, UQVN_N148,
	 UQVN_N149, UQVN_N150, UQVN_N151, UQVN_N152,
	 UQVN_N153, UQVN_N154, UQVN_N155, UQVN_N156,
	 UQVN_N157, UQVN_N158, UQVN_N159, UQVN_N160,
	 UQVN_N161, UQVN_N162, UQVN_N163, UQVN_N164,
	 UQVN_N165, UQVN_N166, UQVN_N167, UQVN_N168,
	 UQVN_N169, UQVN_N170, UQVN_N171, UQVN_N172,
	 UQVN_N173, UQVN_N174, UQVN_N175, UQVN_N176,
	 UQVN_N177, UQVN_N178, UQVN_N179, UQVN_N180,
	 UQVN_N181, UQVN_N182, UQVN_N183, UQVN_N184,
	 UQVN_N185, UQVN_N186, UQVN_N187, UQVN_N188,
	 UQVN_N189, UQVN_N190, UQVN_N191, UQVN_N192,
	 UQVN_N193, UQVN_N194, UQVN_N195, UQVN_N196,
	 UQVN_N197, UQVN_N198, UQVN_N199, UQVN_N200,
	 UQVN_N201, UQVN_N202, UQVN_N203, UQVN_N204,
	 UQVN_N205, UQVN_N206, UQVN_N207, UQVN_N208,
	 UQVN_N209, UQVN_N210, UQVN_N211, UQVN_N212,
	 UQVN_N213, UQVN_N214, UQVN_N215, UQVN_N216,
	 UQVN_N217, UQVN_N218, UQVN_N219, G012,
	 G1214, G345, G678, G911,
	 P1214, P345, P678, P911 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => G012);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B4);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B5);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => A3);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N40, A1 => G012);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => B3, A1 => UQVN_N43);
UQVB_B7 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N3);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N37, A1 => B4, A2 => UQVN_N40);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N41, A1 => B3, A2 => G012);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => A3, A1 => UQVN_N41, A2 => G012);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B4, A1 => UQVN_N40, A2 => UQVN_N43);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N37, A1 => B4, A2 => UQVN_N43);
UQVB_B14 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N8);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A3, A1 => UQVN_N41, A2 => B3);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => A3, A1 => A4, A2 => A5, 
	A3 => B3);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A4, A1 => A5, A2 => B4);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => A3, A1 => A5, A2 => B3, 
	A3 => B4);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A5, A1 => B5);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => A3, A1 => A4, A2 => B3, 
	A3 => B5);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => A4, A1 => B4, A2 => B5);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => A3, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B24 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16, A6 => UQVN_N17);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N37, A1 => UQVN_N40);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N38, A1 => UQVN_N41);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N39, A1 => UQVN_N42);
UQVB_B28 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N20, A1 => UQVN_N18, A2 => UQVN_N19);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => B3);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A4);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A5);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N34);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N41, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N38, A1 => UQVN_N40, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N37, A1 => UQVN_N38, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => B3, A1 => B4, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => A3, A1 => B4, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A4, A1 => B3, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => A3, A1 => A4, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => A3, A1 => B3, A2 => B4, 
	A3 => UQVN_N42);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => A4, A1 => B4, A2 => UQVN_N42);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => A3, A1 => A4, A2 => B3, 
	A3 => UQVN_N42);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N37, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => B5);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N38, A1 => UQVN_N41, A2 => B5);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N37, A1 => UQVN_N38, A2 => UQVN_N40, 
	A3 => B5);
UQVB_B47 : OR12
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N28, A5 => UQVN_N27, A6 => UQVN_N26, 
	A7 => UQVN_N25, A8 => UQVN_N24, A9 => UQVN_N23, A10 => UQVN_N22, 
	A11 => UQVN_N21);
UQVB_B48 : OR3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N33, A1 => UQVN_N35, A2 => UQVN_N36);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N86, A0 => UQVN_N217);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N84, A0 => B10);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N85, A0 => B11);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N80, A0 => A9);
UQVB_B53 : AND2
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N83, A1 => UQVN_N217);
UQVB_B54 : AND2
	PORT MAP (Z0 => UQVN_N45, A0 => B9, A1 => UQVN_N86);
UQVB_B55 : OR2
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N44, A1 => UQVN_N45);
UQVB_B56 : LXOR2
	PORT MAP (Z0 => Z9, A0 => A9, A1 => UQVN_N46);
UQVB_B57 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N80, A1 => B10, A2 => UQVN_N83);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N84, A1 => B9, A2 => UQVN_N217);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N47, A0 => A9, A1 => UQVN_N84, A2 => UQVN_N217);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N49, A0 => B10, A1 => UQVN_N83, A2 => UQVN_N86);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N80, A1 => B10, A2 => UQVN_N86);
UQVB_B62 : OR6
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N50, A1 => UQVN_N49, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N52, A5 => UQVN_N51);
UQVB_B63 : LXOR2
	PORT MAP (Z0 => Z10, A0 => A10, A1 => UQVN_N53);
UQVB_B64 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => A9, A1 => UQVN_N84, A2 => B9);
UQVB_B65 : AND4
	PORT MAP (Z0 => UQVN_N57, A0 => A9, A1 => A10, A2 => A11, 
	A3 => B9);
UQVB_B66 : AND3
	PORT MAP (Z0 => UQVN_N56, A0 => A10, A1 => A11, A2 => B10);
UQVB_B67 : AND4
	PORT MAP (Z0 => UQVN_N55, A0 => A9, A1 => A11, A2 => B9, 
	A3 => B10);
UQVB_B68 : AND2
	PORT MAP (Z0 => UQVN_N54, A0 => A11, A1 => B11);
UQVB_B69 : AND4
	PORT MAP (Z0 => UQVN_N58, A0 => A9, A1 => A10, A2 => B9, 
	A3 => B11);
UQVB_B70 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => A10, A1 => B10, A2 => B11);
UQVB_B71 : AND4
	PORT MAP (Z0 => UQVN_N60, A0 => A9, A1 => B9, A2 => B10, 
	A3 => B11);
UQVB_B72 : OR7
	PORT MAP (Z0 => G911, A0 => UQVN_N57, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N58, A5 => UQVN_N59, A6 => UQVN_N60);
UQVB_B73 : AND2
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N80, A1 => UQVN_N83);
UQVB_B74 : AND2
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N81, A1 => UQVN_N84);
UQVB_B75 : AND2
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N82, A1 => UQVN_N85);
UQVB_B76 : NOR3
	PORT MAP (ZN0 => P911, A0 => UQVN_N63, A1 => UQVN_N61, A2 => UQVN_N62);
UQVB_B77 : INV
	PORT MAP (ZN0 => UQVN_N83, A0 => B9);
UQVB_B78 : INV
	PORT MAP (ZN0 => UQVN_N81, A0 => A10);
UQVB_B79 : INV
	PORT MAP (ZN0 => UQVN_N82, A0 => A11);
UQVB_B80 : LXOR2
	PORT MAP (Z0 => Z11, A0 => A11, A1 => UQVN_N77);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N83, A1 => UQVN_N84, A2 => B11, 
	A3 => UQVN_N86);
UQVB_B82 : AND4
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N80, A1 => UQVN_N84, A2 => B11, 
	A3 => UQVN_N86);
UQVB_B83 : AND4
	PORT MAP (Z0 => UQVN_N75, A0 => UQVN_N81, A1 => UQVN_N83, A2 => B11, 
	A3 => UQVN_N86);
UQVB_B84 : AND4
	PORT MAP (Z0 => UQVN_N74, A0 => UQVN_N80, A1 => UQVN_N81, A2 => B11, 
	A3 => UQVN_N86);
UQVB_B85 : AND4
	PORT MAP (Z0 => UQVN_N73, A0 => B9, A1 => B10, A2 => UQVN_N85, 
	A3 => UQVN_N217);
UQVB_B86 : AND4
	PORT MAP (Z0 => UQVN_N72, A0 => A9, A1 => B10, A2 => UQVN_N85, 
	A3 => UQVN_N217);
UQVB_B87 : AND4
	PORT MAP (Z0 => UQVN_N71, A0 => A10, A1 => B9, A2 => UQVN_N85, 
	A3 => UQVN_N217);
UQVB_B88 : AND4
	PORT MAP (Z0 => UQVN_N70, A0 => A9, A1 => A10, A2 => UQVN_N85, 
	A3 => UQVN_N217);
UQVB_B89 : AND4
	PORT MAP (Z0 => UQVN_N69, A0 => A9, A1 => B9, A2 => B10, 
	A3 => UQVN_N85);
UQVB_B90 : AND3
	PORT MAP (Z0 => UQVN_N68, A0 => A10, A1 => B10, A2 => UQVN_N85);
UQVB_B91 : AND4
	PORT MAP (Z0 => UQVN_N67, A0 => A9, A1 => A10, A2 => B9, 
	A3 => UQVN_N85);
UQVB_B92 : AND4
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N80, A1 => UQVN_N83, A2 => UQVN_N84, 
	A3 => B11);
UQVB_B93 : AND3
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N81, A1 => UQVN_N84, A2 => B11);
UQVB_B94 : AND4
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N80, A1 => UQVN_N81, A2 => UQVN_N83, 
	A3 => B11);
UQVB_B95 : OR12
	PORT MAP (Z0 => UQVN_N79, A0 => UQVN_N75, A1 => UQVN_N74, A2 => UQVN_N73, 
	A3 => UQVN_N72, A4 => UQVN_N71, A5 => UQVN_N70, A6 => UQVN_N69, 
	A7 => UQVN_N68, A8 => UQVN_N67, A9 => UQVN_N66, A10 => UQVN_N65, 
	A11 => UQVN_N64);
UQVB_B96 : OR3
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N76, A1 => UQVN_N78, A2 => UQVN_N79);
UQVB_B97 : INV
	PORT MAP (ZN0 => UQVN_N129, A0 => UQVN_N218);
UQVB_B98 : INV
	PORT MAP (ZN0 => UQVN_N127, A0 => B13);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N128, A0 => B14);
UQVB_B100 : INV
	PORT MAP (ZN0 => UQVN_N123, A0 => A12);
UQVB_B101 : AND2
	PORT MAP (Z0 => UQVN_N87, A0 => UQVN_N126, A1 => UQVN_N218);
UQVB_B102 : AND2
	PORT MAP (Z0 => UQVN_N88, A0 => B12, A1 => UQVN_N129);
UQVB_B103 : OR2
	PORT MAP (Z0 => UQVN_N89, A0 => UQVN_N87, A1 => UQVN_N88);
UQVB_B104 : LXOR2
	PORT MAP (Z0 => Z12, A0 => A12, A1 => UQVN_N89);
UQVB_B105 : AND3
	PORT MAP (Z0 => UQVN_N95, A0 => UQVN_N123, A1 => B13, A2 => UQVN_N126);
UQVB_B106 : AND3
	PORT MAP (Z0 => UQVN_N91, A0 => UQVN_N127, A1 => B12, A2 => UQVN_N218);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N90, A0 => A12, A1 => UQVN_N127, A2 => UQVN_N218);
UQVB_B108 : AND3
	PORT MAP (Z0 => UQVN_N92, A0 => B13, A1 => UQVN_N126, A2 => UQVN_N129);
UQVB_B109 : AND3
	PORT MAP (Z0 => UQVN_N93, A0 => UQVN_N123, A1 => B13, A2 => UQVN_N129);
UQVB_B110 : OR6
	PORT MAP (Z0 => UQVN_N96, A0 => UQVN_N93, A1 => UQVN_N92, A2 => UQVN_N90, 
	A3 => UQVN_N91, A4 => UQVN_N95, A5 => UQVN_N94);
UQVB_B111 : LXOR2
	PORT MAP (Z0 => Z13, A0 => A13, A1 => UQVN_N96);
UQVB_B112 : AND3
	PORT MAP (Z0 => UQVN_N94, A0 => A12, A1 => UQVN_N127, A2 => B12);
UQVB_B113 : AND4
	PORT MAP (Z0 => UQVN_N100, A0 => A12, A1 => A13, A2 => A14, 
	A3 => B12);
UQVB_B114 : AND3
	PORT MAP (Z0 => UQVN_N99, A0 => A13, A1 => A14, A2 => B13);
UQVB_B115 : AND4
	PORT MAP (Z0 => UQVN_N98, A0 => A12, A1 => A14, A2 => B12, 
	A3 => B13);
UQVB_B116 : AND2
	PORT MAP (Z0 => UQVN_N97, A0 => A14, A1 => B14);
UQVB_B117 : AND4
	PORT MAP (Z0 => UQVN_N101, A0 => A12, A1 => A13, A2 => B12, 
	A3 => B14);
UQVB_B118 : AND3
	PORT MAP (Z0 => UQVN_N102, A0 => A13, A1 => B13, A2 => B14);
UQVB_B119 : AND4
	PORT MAP (Z0 => UQVN_N103, A0 => A12, A1 => B12, A2 => B13, 
	A3 => B14);
UQVB_B120 : OR7
	PORT MAP (Z0 => G1214, A0 => UQVN_N100, A1 => UQVN_N99, A2 => UQVN_N98, 
	A3 => UQVN_N97, A4 => UQVN_N101, A5 => UQVN_N102, A6 => UQVN_N103);
UQVB_B121 : AND2
	PORT MAP (Z0 => UQVN_N106, A0 => UQVN_N123, A1 => UQVN_N126);
UQVB_B122 : AND2
	PORT MAP (Z0 => UQVN_N104, A0 => UQVN_N124, A1 => UQVN_N127);
UQVB_B123 : AND2
	PORT MAP (Z0 => UQVN_N105, A0 => UQVN_N125, A1 => UQVN_N128);
UQVB_B124 : NOR3
	PORT MAP (ZN0 => P1214, A0 => UQVN_N106, A1 => UQVN_N104, A2 => UQVN_N105);
UQVB_B125 : INV
	PORT MAP (ZN0 => UQVN_N126, A0 => B12);
UQVB_B126 : INV
	PORT MAP (ZN0 => UQVN_N124, A0 => A13);
UQVB_B127 : INV
	PORT MAP (ZN0 => UQVN_N125, A0 => A14);
UQVB_B128 : LXOR2
	PORT MAP (Z0 => Z14, A0 => A14, A1 => UQVN_N120);
UQVB_B129 : AND4
	PORT MAP (Z0 => UQVN_N119, A0 => UQVN_N126, A1 => UQVN_N127, A2 => B14, 
	A3 => UQVN_N129);
UQVB_B130 : AND4
	PORT MAP (Z0 => UQVN_N121, A0 => UQVN_N123, A1 => UQVN_N127, A2 => B14, 
	A3 => UQVN_N129);
UQVB_B131 : AND4
	PORT MAP (Z0 => UQVN_N118, A0 => UQVN_N124, A1 => UQVN_N126, A2 => B14, 
	A3 => UQVN_N129);
UQVB_B132 : AND4
	PORT MAP (Z0 => UQVN_N117, A0 => UQVN_N123, A1 => UQVN_N124, A2 => B14, 
	A3 => UQVN_N129);
UQVB_B133 : AND4
	PORT MAP (Z0 => UQVN_N116, A0 => B12, A1 => B13, A2 => UQVN_N128, 
	A3 => UQVN_N218);
UQVB_B134 : AND4
	PORT MAP (Z0 => UQVN_N115, A0 => A12, A1 => B13, A2 => UQVN_N128, 
	A3 => UQVN_N218);
UQVB_B135 : AND4
	PORT MAP (Z0 => UQVN_N114, A0 => A13, A1 => B12, A2 => UQVN_N128, 
	A3 => UQVN_N218);
UQVB_B136 : AND4
	PORT MAP (Z0 => UQVN_N113, A0 => A12, A1 => A13, A2 => UQVN_N128, 
	A3 => UQVN_N218);
UQVB_B137 : AND4
	PORT MAP (Z0 => UQVN_N112, A0 => A12, A1 => B12, A2 => B13, 
	A3 => UQVN_N128);
UQVB_B138 : AND3
	PORT MAP (Z0 => UQVN_N111, A0 => A13, A1 => B13, A2 => UQVN_N128);
UQVB_B139 : AND4
	PORT MAP (Z0 => UQVN_N110, A0 => A12, A1 => A13, A2 => B12, 
	A3 => UQVN_N128);
UQVB_B140 : AND4
	PORT MAP (Z0 => UQVN_N109, A0 => UQVN_N123, A1 => UQVN_N126, A2 => UQVN_N127, 
	A3 => B14);
UQVB_B141 : AND3
	PORT MAP (Z0 => UQVN_N108, A0 => UQVN_N124, A1 => UQVN_N127, A2 => B14);
UQVB_B142 : AND4
	PORT MAP (Z0 => UQVN_N107, A0 => UQVN_N123, A1 => UQVN_N124, A2 => UQVN_N126, 
	A3 => B14);
UQVB_B143 : OR12
	PORT MAP (Z0 => UQVN_N122, A0 => UQVN_N118, A1 => UQVN_N117, A2 => UQVN_N116, 
	A3 => UQVN_N115, A4 => UQVN_N114, A5 => UQVN_N113, A6 => UQVN_N112, 
	A7 => UQVN_N111, A8 => UQVN_N110, A9 => UQVN_N109, A10 => UQVN_N108, 
	A11 => UQVN_N107);
UQVB_B144 : OR3
	PORT MAP (Z0 => UQVN_N120, A0 => UQVN_N119, A1 => UQVN_N121, A2 => UQVN_N122);
UQVB_B145 : AND2
	PORT MAP (Z0 => UQVN_N130, A0 => P345, A1 => G012);
UQVB_B146 : OR2
	PORT MAP (Z0 => UQVN_N216, A0 => G345, A1 => UQVN_N130);
UQVB_B147 : INV
	PORT MAP (ZN0 => UQVN_N173, A0 => UQVN_N216);
UQVB_B148 : INV
	PORT MAP (ZN0 => UQVN_N171, A0 => B7);
UQVB_B149 : INV
	PORT MAP (ZN0 => UQVN_N172, A0 => B8);
UQVB_B150 : INV
	PORT MAP (ZN0 => UQVN_N167, A0 => A6);
UQVB_B151 : AND2
	PORT MAP (Z0 => UQVN_N131, A0 => UQVN_N170, A1 => UQVN_N216);
UQVB_B152 : AND2
	PORT MAP (Z0 => UQVN_N132, A0 => B6, A1 => UQVN_N173);
UQVB_B153 : OR2
	PORT MAP (Z0 => UQVN_N133, A0 => UQVN_N131, A1 => UQVN_N132);
UQVB_B154 : LXOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N133);
UQVB_B155 : AND3
	PORT MAP (Z0 => UQVN_N139, A0 => UQVN_N167, A1 => B7, A2 => UQVN_N170);
UQVB_B156 : AND3
	PORT MAP (Z0 => UQVN_N135, A0 => UQVN_N171, A1 => B6, A2 => UQVN_N216);
UQVB_B157 : AND3
	PORT MAP (Z0 => UQVN_N134, A0 => A6, A1 => UQVN_N171, A2 => UQVN_N216);
UQVB_B158 : AND3
	PORT MAP (Z0 => UQVN_N136, A0 => B7, A1 => UQVN_N170, A2 => UQVN_N173);
UQVB_B159 : AND3
	PORT MAP (Z0 => UQVN_N137, A0 => UQVN_N167, A1 => B7, A2 => UQVN_N173);
UQVB_B160 : OR6
	PORT MAP (Z0 => UQVN_N140, A0 => UQVN_N137, A1 => UQVN_N136, A2 => UQVN_N134, 
	A3 => UQVN_N135, A4 => UQVN_N139, A5 => UQVN_N138);
UQVB_B161 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N140);
UQVB_B162 : AND3
	PORT MAP (Z0 => UQVN_N138, A0 => A6, A1 => UQVN_N171, A2 => B6);
UQVB_B163 : AND4
	PORT MAP (Z0 => UQVN_N144, A0 => A6, A1 => A7, A2 => A8, 
	A3 => B6);
UQVB_B164 : AND3
	PORT MAP (Z0 => UQVN_N143, A0 => A7, A1 => A8, A2 => B7);
UQVB_B165 : AND4
	PORT MAP (Z0 => UQVN_N142, A0 => A6, A1 => A8, A2 => B6, 
	A3 => B7);
UQVB_B166 : AND2
	PORT MAP (Z0 => UQVN_N141, A0 => A8, A1 => B8);
UQVB_B167 : AND4
	PORT MAP (Z0 => UQVN_N145, A0 => A6, A1 => A7, A2 => B6, 
	A3 => B8);
UQVB_B168 : AND3
	PORT MAP (Z0 => UQVN_N146, A0 => A7, A1 => B7, A2 => B8);
UQVB_B169 : AND4
	PORT MAP (Z0 => UQVN_N147, A0 => A6, A1 => B6, A2 => B7, 
	A3 => B8);
UQVB_B170 : OR7
	PORT MAP (Z0 => G678, A0 => UQVN_N144, A1 => UQVN_N143, A2 => UQVN_N142, 
	A3 => UQVN_N141, A4 => UQVN_N145, A5 => UQVN_N146, A6 => UQVN_N147);
UQVB_B171 : AND2
	PORT MAP (Z0 => UQVN_N150, A0 => UQVN_N167, A1 => UQVN_N170);
UQVB_B172 : AND2
	PORT MAP (Z0 => UQVN_N148, A0 => UQVN_N168, A1 => UQVN_N171);
UQVB_B173 : AND2
	PORT MAP (Z0 => UQVN_N149, A0 => UQVN_N169, A1 => UQVN_N172);
UQVB_B174 : NOR3
	PORT MAP (ZN0 => P678, A0 => UQVN_N150, A1 => UQVN_N148, A2 => UQVN_N149);
UQVB_B175 : INV
	PORT MAP (ZN0 => UQVN_N170, A0 => B6);
UQVB_B176 : INV
	PORT MAP (ZN0 => UQVN_N168, A0 => A7);
UQVB_B177 : INV
	PORT MAP (ZN0 => UQVN_N169, A0 => A8);
UQVB_B178 : LXOR2
	PORT MAP (Z0 => Z8, A0 => A8, A1 => UQVN_N164);
UQVB_B179 : AND4
	PORT MAP (Z0 => UQVN_N163, A0 => UQVN_N170, A1 => UQVN_N171, A2 => B8, 
	A3 => UQVN_N173);
UQVB_B180 : AND4
	PORT MAP (Z0 => UQVN_N165, A0 => UQVN_N167, A1 => UQVN_N171, A2 => B8, 
	A3 => UQVN_N173);
UQVB_B181 : AND4
	PORT MAP (Z0 => UQVN_N162, A0 => UQVN_N168, A1 => UQVN_N170, A2 => B8, 
	A3 => UQVN_N173);
UQVB_B182 : AND4
	PORT MAP (Z0 => UQVN_N161, A0 => UQVN_N167, A1 => UQVN_N168, A2 => B8, 
	A3 => UQVN_N173);
UQVB_B183 : AND4
	PORT MAP (Z0 => UQVN_N160, A0 => B6, A1 => B7, A2 => UQVN_N172, 
	A3 => UQVN_N216);
UQVB_B184 : AND4
	PORT MAP (Z0 => UQVN_N159, A0 => A6, A1 => B7, A2 => UQVN_N172, 
	A3 => UQVN_N216);
UQVB_B185 : AND4
	PORT MAP (Z0 => UQVN_N158, A0 => A7, A1 => B6, A2 => UQVN_N172, 
	A3 => UQVN_N216);
UQVB_B186 : AND4
	PORT MAP (Z0 => UQVN_N157, A0 => A6, A1 => A7, A2 => UQVN_N172, 
	A3 => UQVN_N216);
UQVB_B187 : AND4
	PORT MAP (Z0 => UQVN_N156, A0 => A6, A1 => B6, A2 => B7, 
	A3 => UQVN_N172);
UQVB_B188 : AND3
	PORT MAP (Z0 => UQVN_N155, A0 => A7, A1 => B7, A2 => UQVN_N172);
UQVB_B189 : AND4
	PORT MAP (Z0 => UQVN_N154, A0 => A6, A1 => A7, A2 => B6, 
	A3 => UQVN_N172);
UQVB_B190 : AND4
	PORT MAP (Z0 => UQVN_N153, A0 => UQVN_N167, A1 => UQVN_N170, A2 => UQVN_N171, 
	A3 => B8);
UQVB_B191 : AND3
	PORT MAP (Z0 => UQVN_N152, A0 => UQVN_N168, A1 => UQVN_N171, A2 => B8);
UQVB_B192 : AND4
	PORT MAP (Z0 => UQVN_N151, A0 => UQVN_N167, A1 => UQVN_N168, A2 => UQVN_N170, 
	A3 => B8);
UQVB_B193 : OR12
	PORT MAP (Z0 => UQVN_N166, A0 => UQVN_N162, A1 => UQVN_N161, A2 => UQVN_N160, 
	A3 => UQVN_N159, A4 => UQVN_N158, A5 => UQVN_N157, A6 => UQVN_N156, 
	A7 => UQVN_N155, A8 => UQVN_N154, A9 => UQVN_N153, A10 => UQVN_N152, 
	A11 => UQVN_N151);
UQVB_B194 : OR3
	PORT MAP (Z0 => UQVN_N164, A0 => UQVN_N163, A1 => UQVN_N165, A2 => UQVN_N166);
UQVB_B195 : OR3
	PORT MAP (Z0 => UQVN_N217, A0 => G678, A1 => UQVN_N174, A2 => UQVN_N175);
UQVB_B196 : AND3
	PORT MAP (Z0 => UQVN_N175, A0 => P678, A1 => P345, A2 => G012);
UQVB_B197 : AND2
	PORT MAP (Z0 => UQVN_N174, A0 => P678, A1 => G345);
UQVB_B198 : OR4
	PORT MAP (Z0 => UQVN_N218, A0 => G911, A1 => UQVN_N176, A2 => UQVN_N177, 
	A3 => UQVN_N178);
UQVB_B199 : AND2
	PORT MAP (Z0 => UQVN_N176, A0 => P911, A1 => G678);
UQVB_B200 : AND3
	PORT MAP (Z0 => UQVN_N177, A0 => P911, A1 => P678, A2 => G345);
UQVB_B201 : AND4
	PORT MAP (Z0 => UQVN_N178, A0 => P911, A1 => P678, A2 => P345, 
	A3 => G012);
UQVB_B202 : OR5
	PORT MAP (Z0 => UQVN_N219, A0 => G1214, A1 => UQVN_N179, A2 => UQVN_N180, 
	A3 => UQVN_N181, A4 => UQVN_N182);
UQVB_B203 : AND2
	PORT MAP (Z0 => UQVN_N179, A0 => P1214, A1 => G911);
UQVB_B204 : AND3
	PORT MAP (Z0 => UQVN_N180, A0 => P1214, A1 => P911, A2 => G678);
UQVB_B205 : AND4
	PORT MAP (Z0 => UQVN_N181, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => G345);
UQVB_B206 : AND5
	PORT MAP (Z0 => UQVN_N182, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => P345, A4 => G012);
UQVB_B207 : INV
	PORT MAP (ZN0 => UQVN_N206, A0 => B1);
UQVB_B208 : INV
	PORT MAP (ZN0 => UQVN_N203, A0 => A0);
UQVB_B209 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B210 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N186);
UQVB_B211 : AND3
	PORT MAP (Z0 => UQVN_N185, A0 => A0, A1 => UQVN_N206, A2 => B0);
UQVB_B212 : AND4
	PORT MAP (Z0 => UQVN_N190, A0 => A0, A1 => A1, A2 => A2, 
	A3 => B0);
UQVB_B213 : AND3
	PORT MAP (Z0 => UQVN_N189, A0 => A1, A1 => A2, A2 => B1);
UQVB_B214 : AND4
	PORT MAP (Z0 => UQVN_N188, A0 => A0, A1 => A2, A2 => B0, 
	A3 => B1);
UQVB_B215 : AND2
	PORT MAP (Z0 => UQVN_N187, A0 => A2, A1 => B2);
UQVB_B216 : AND4
	PORT MAP (Z0 => UQVN_N191, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B2);
UQVB_B217 : AND3
	PORT MAP (Z0 => UQVN_N192, A0 => A1, A1 => B1, A2 => B2);
UQVB_B218 : AND4
	PORT MAP (Z0 => UQVN_N193, A0 => A0, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B219 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N190, A1 => UQVN_N189, A2 => UQVN_N188, 
	A3 => UQVN_N187, A4 => UQVN_N191, A5 => UQVN_N192, A6 => UQVN_N193);
UQVB_B220 : INV
	PORT MAP (ZN0 => UQVN_N205, A0 => B0);
UQVB_B221 : INV
	PORT MAP (ZN0 => UQVN_N204, A0 => A1);
UQVB_B222 : AND2
	PORT MAP (Z0 => UQVN_N184, A0 => UQVN_N203, A1 => B1);
UQVB_B223 : AND2
	PORT MAP (Z0 => UQVN_N183, A0 => B1, A1 => UQVN_N205);
UQVB_B224 : OR3
	PORT MAP (Z0 => UQVN_N186, A0 => UQVN_N184, A1 => UQVN_N183, A2 => UQVN_N185);
UQVB_B225 : INV
	PORT MAP (ZN0 => UQVN_N207, A0 => B2);
UQVB_B226 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N198);
UQVB_B227 : AND4
	PORT MAP (Z0 => UQVN_N197, A0 => A0, A1 => B0, A2 => B1, 
	A3 => UQVN_N207);
UQVB_B228 : AND3
	PORT MAP (Z0 => UQVN_N196, A0 => A1, A1 => B1, A2 => UQVN_N207);
UQVB_B229 : AND4
	PORT MAP (Z0 => UQVN_N195, A0 => A0, A1 => A1, A2 => B0, 
	A3 => UQVN_N207);
UQVB_B230 : AND3
	PORT MAP (Z0 => UQVN_N194, A0 => UQVN_N204, A1 => UQVN_N206, A2 => B2);
UQVB_B231 : AND3
	PORT MAP (Z0 => UQVN_N202, A0 => UQVN_N205, A1 => UQVN_N206, A2 => B2);
UQVB_B232 : AND3
	PORT MAP (Z0 => UQVN_N201, A0 => UQVN_N203, A1 => UQVN_N206, A2 => B2);
UQVB_B233 : AND3
	PORT MAP (Z0 => UQVN_N200, A0 => UQVN_N204, A1 => UQVN_N205, A2 => B2);
UQVB_B234 : AND3
	PORT MAP (Z0 => UQVN_N199, A0 => UQVN_N203, A1 => UQVN_N204, A2 => B2);
UQVB_B235 : OR8
	PORT MAP (Z0 => UQVN_N198, A0 => UQVN_N202, A1 => UQVN_N201, A2 => UQVN_N200, 
	A3 => UQVN_N199, A4 => UQVN_N197, A5 => UQVN_N196, A6 => UQVN_N195, 
	A7 => UQVN_N194);
UQVB_B236 : AND2
	PORT MAP (Z0 => UQVN_N209, A0 => UQVN_N215, A1 => UQVN_N219);
UQVB_B237 : AND2
	PORT MAP (Z0 => UQVN_N210, A0 => B15, A1 => UQVN_N208);
UQVB_B238 : OR2
	PORT MAP (Z0 => UQVN_N211, A0 => UQVN_N210, A1 => UQVN_N209);
UQVB_B239 : XOR2
	PORT MAP (Z0 => Z15, A0 => A15, A1 => UQVN_N211);
UQVB_B240 : INV
	PORT MAP (ZN0 => UQVN_N215, A0 => B15);
UQVB_B241 : INV
	PORT MAP (ZN0 => UQVN_N208, A0 => UQVN_N219);
UQVB_B242 : AND2
	PORT MAP (Z0 => UQVN_N212, A0 => UQVN_N219, A1 => B15);
UQVB_B243 : AND2
	PORT MAP (Z0 => UQVN_N213, A0 => UQVN_N219, A1 => A15);
UQVB_B244 : AND2
	PORT MAP (Z0 => UQVN_N214, A0 => B15, A1 => A15);
UQVB_B245 : OR3
	PORT MAP (Z0 => CO, A0 => UQVN_N212, A1 => UQVN_N213, A2 => UQVN_N214);
END lattice_arch;
-- VHDL netlist for ADDH2
-- Date: 15.5.95 13.44.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDH2;


ARCHITECTURE lattice_arch OF ADDH2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N12, A1 => B0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N14);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => A1, A1 => A0, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => B1, A2 => B0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => A1, A1 => B1);
UQVB_B6 : OR3
	PORT MAP (Z0 => CO, A0 => UQVN_N3, A1 => UQVN_N5, A2 => UQVN_N4);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => B0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => B1);
UQVB_B10 : OR6
	PORT MAP (Z0 => Z1, A0 => UQVN_N6, A1 => UQVN_N8, A2 => UQVN_N7, 
	A3 => UQVN_N9, A4 => UQVN_N10, A5 => UQVN_N11);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N13, A1 => B1, A2 => UQVN_N12);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N13, A1 => B1, A2 => UQVN_N14);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N15, A2 => UQVN_N12);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => A1, A1 => UQVN_N15, A2 => UQVN_N14);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N13, A1 => UQVN_N15, A2 => A0, 
	A3 => B0);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A1, A1 => B1, A2 => A0, 
	A3 => B0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => A0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => A1);
END lattice_arch;
-- VHDL netlist for ADDH3
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH3 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDH3;


ARCHITECTURE lattice_arch OF ADDH3 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => B1);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => A0);
UQVB_B3 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B4 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N4);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => A0, A1 => UQVN_N24, A2 => B0);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => A1, A2 => A2, 
	A3 => B0);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => A2, A2 => B1);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => A0, A1 => A2, A2 => B0, 
	A3 => B1);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => A2, A1 => B2);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B2);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => A1, A1 => B1, A2 => B2);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A0, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B13 : OR7
	PORT MAP (Z0 => CO, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N10, A6 => UQVN_N11);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => B0);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => A1);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N21, A1 => B1);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => B1, A1 => UQVN_N23);
UQVB_B18 : OR3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => B2);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N16);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => A0, A1 => B0, A2 => B1, 
	A3 => UQVN_N25);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => A1, A1 => B1, A2 => UQVN_N25);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => A0, A1 => A1, A2 => B0, 
	A3 => UQVN_N25);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N22, A1 => UQVN_N24, A2 => B2);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N23, A1 => UQVN_N24, A2 => B2);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N21, A1 => UQVN_N24, A2 => B2);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N22, A1 => UQVN_N23, A2 => B2);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N21, A1 => UQVN_N22, A2 => B2);
UQVB_B29 : OR8
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N18, 
	A3 => UQVN_N17, A4 => UQVN_N15, A5 => UQVN_N14, A6 => UQVN_N13, 
	A7 => UQVN_N12);
END lattice_arch;
-- VHDL netlist for ADDH4
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDH4;


ARCHITECTURE lattice_arch OF ADDH4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N12, A1 => B0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N14);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => A1, A1 => A0, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => B1, A2 => B0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => A1, A1 => B1);
UQVB_B6 : OR3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N3, A1 => UQVN_N5, A2 => UQVN_N4);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => B0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => B1);
UQVB_B10 : OR6
	PORT MAP (Z0 => Z1, A0 => UQVN_N6, A1 => UQVN_N8, A2 => UQVN_N7, 
	A3 => UQVN_N9, A4 => UQVN_N10, A5 => UQVN_N11);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N13, A1 => B1, A2 => UQVN_N12);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N13, A1 => B1, A2 => UQVN_N14);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N15, A2 => UQVN_N12);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => A1, A1 => UQVN_N15, A2 => UQVN_N14);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N13, A1 => UQVN_N15, A2 => A0, 
	A3 => B0);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A1, A1 => B1, A2 => A0, 
	A3 => B0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => A0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => A1);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => UQVN_N37);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N37, A1 => A3, A2 => A2);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N37, A1 => A3, A2 => B2);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N37, A1 => A2, A2 => B3);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N37, A1 => B3, A2 => B2);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => A3, A1 => A2, A2 => B2);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => A2, A1 => B3, A2 => B2);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => A3, A1 => B3);
UQVB_B27 : OR7
	PORT MAP (Z0 => CO, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N16, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => UQVN_N22, A6 => UQVN_N21);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N33, A1 => B3, A2 => UQVN_N36);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => B3, A1 => UQVN_N34, A2 => UQVN_N36);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => A2, A1 => UQVN_N35, A2 => UQVN_N37);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N35, A1 => B2, A2 => UQVN_N37);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N33, A1 => B3, A2 => UQVN_N34);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => A2, A1 => UQVN_N35, A2 => B2);
UQVB_B34 : OR6
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N23, A1 => UQVN_N24, A2 => UQVN_N25, 
	A3 => UQVN_N26, A4 => UQVN_N27, A5 => UQVN_N28);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N29);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => B2);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => B3);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => A2);
UQVB_B39 : XOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N30);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N37, A1 => UQVN_N34);
UQVB_B41 : OR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N31, A1 => UQVN_N32);
UQVB_B42 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => B2);
END lattice_arch;
-- VHDL netlist for ADDH8
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        CO : OUT std_logic
    );
END ADDH8;


ARCHITECTURE lattice_arch OF ADDH8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, G1, G2, G3,
	 G4, G5, G6, G7,
	 P1, P2, P3, P4,
	 P5, P6, P7 : std_logic;


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : XOR2
	PORT MAP (Z0 => P7, A0 => A7, A1 => B7);
UQVB_B2 : XOR2
	PORT MAP (Z0 => P6, A0 => A6, A1 => B6);
UQVB_B3 : XOR2
	PORT MAP (Z0 => P5, A0 => A5, A1 => B5);
UQVB_B4 : XOR2
	PORT MAP (Z0 => P4, A0 => A4, A1 => B4);
UQVB_B5 : XOR2
	PORT MAP (Z0 => P3, A0 => A3, A1 => B3);
UQVB_B6 : XOR2
	PORT MAP (Z0 => P2, A0 => A2, A1 => B2);
UQVB_B7 : XOR2
	PORT MAP (Z0 => P1, A0 => A1, A1 => B1);
UQVB_B8 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B9 : AND2
	PORT MAP (Z0 => G7, A0 => A7, A1 => B7);
UQVB_B10 : AND2
	PORT MAP (Z0 => G6, A0 => A6, A1 => B6);
UQVB_B11 : AND2
	PORT MAP (Z0 => G5, A0 => A5, A1 => B5);
UQVB_B12 : AND2
	PORT MAP (Z0 => G4, A0 => A4, A1 => B4);
UQVB_B13 : AND2
	PORT MAP (Z0 => G3, A0 => A3, A1 => B3);
UQVB_B14 : AND2
	PORT MAP (Z0 => G2, A0 => A2, A1 => B2);
UQVB_B15 : AND2
	PORT MAP (Z0 => G1, A0 => A1, A1 => B1);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => B0);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => Z1, A0 => P1, A1 => UQVN_N1);
UQVB_B18 : AND9
	PORT MAP (Z0 => UQVN_N13, A0 => A0, A1 => B0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4, A6 => P5, 
	A7 => P6, A8 => P7);
UQVB_B19 : OR5
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => G4);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N6, A1 => P5);
UQVB_B21 : AND7
	PORT MAP (Z0 => UQVN_N12, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4, A4 => P5, A5 => P6, A6 => P7);
UQVB_B22 : OR4
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N15, A1 => UQVN_N18, A2 => UQVN_N17, 
	A3 => G7);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => B0, A2 => P1);
UQVB_B24 : OR2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N8, A1 => G1);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N7, A1 => P2);
UQVB_B26 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N13, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => UQVN_N16);
UQVB_B27 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N11, A1 => UQVN_N9, A2 => G2);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => G1, A1 => P2);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N10, A1 => P3);
UQVB_B30 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A0, A1 => B0, A2 => P1, 
	A3 => P2);
UQVB_B31 : AND6
	PORT MAP (Z0 => UQVN_N14, A0 => G2, A1 => P3, A2 => P4, 
	A3 => P5, A4 => P6, A5 => P7);
UQVB_B32 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => G3, A1 => P4, A2 => P5, 
	A3 => P6, A4 => P7);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => G6, A1 => P7);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => G5, A1 => P6, A2 => P7);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => G4, A1 => P5, A2 => P6, 
	A3 => P7);
UQVB_B36 : OR2
	PORT MAP (Z0 => CO, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B37 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => A0, A1 => B0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4);
UQVB_B39 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => G2, A1 => P3, A2 => P4);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => G3, A1 => P4);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => G3, A1 => P4, A2 => P5);
UQVB_B42 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => G2, A1 => P3, A2 => P4, 
	A3 => P5);
UQVB_B43 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4, A4 => P5);
UQVB_B44 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => G4, A1 => P5);
UQVB_B45 : OR3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N24, A1 => UQVN_N23, A2 => G5);
UQVB_B46 : OR3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N28, A1 => UQVN_N22, A2 => UQVN_N25);
UQVB_B47 : OR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N27, A1 => UQVN_N26);
UQVB_B48 : LXOR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N21, A1 => P6);
UQVB_B49 : AND7
	PORT MAP (Z0 => UQVN_N28, A0 => A0, A1 => B0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4, A6 => P5);
UQVB_B50 : AND5
	PORT MAP (Z0 => UQVN_N32, A0 => A0, A1 => B0, A2 => P1, 
	A3 => P2, A4 => P3);
UQVB_B51 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => G1, A1 => P2, A2 => P3);
UQVB_B52 : AND2
	PORT MAP (Z0 => UQVN_N30, A0 => G2, A1 => P3);
UQVB_B53 : OR4
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N32, A1 => UQVN_N29, A2 => UQVN_N30, 
	A3 => G3);
UQVB_B54 : LXOR2
	PORT MAP (Z0 => Z4, A0 => UQVN_N31, A1 => P4);
UQVB_B55 : OR2
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N34, A1 => UQVN_N33);
UQVB_B56 : AND2
	PORT MAP (Z0 => UQVN_N40, A0 => G5, A1 => P6);
UQVB_B57 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => G4, A1 => P5, A2 => P6);
UQVB_B58 : AND4
	PORT MAP (Z0 => UQVN_N39, A0 => G3, A1 => P4, A2 => P5, 
	A3 => P6);
UQVB_B59 : AND5
	PORT MAP (Z0 => UQVN_N37, A0 => G2, A1 => P3, A2 => P4, 
	A3 => P5, A4 => P6);
UQVB_B60 : AND6
	PORT MAP (Z0 => UQVN_N35, A0 => G1, A1 => P2, A2 => P3, 
	A3 => P4, A4 => P5, A5 => P6);
UQVB_B61 : AND8
	PORT MAP (Z0 => UQVN_N36, A0 => A0, A1 => B0, A2 => P1, 
	A3 => P2, A4 => P3, A5 => P4, A6 => P5, 
	A7 => P6);
UQVB_B62 : OR4
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N36, A1 => UQVN_N35, A2 => UQVN_N37, 
	A3 => UQVN_N39);
UQVB_B63 : OR3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N38, A1 => UQVN_N40, A2 => G6);
UQVB_B64 : LXOR2
	PORT MAP (Z0 => Z7, A0 => UQVN_N41, A1 => P7);
END lattice_arch;
-- VHDL netlist for ADDH8A
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ADDH8A IS 
    PORT (
        B7 : IN std_logic;
        B6 : IN std_logic;
        B5 : IN std_logic;
        B4 : IN std_logic;
        B3 : IN std_logic;
        B2 : IN std_logic;
        B1 : IN std_logic;
        B0 : IN std_logic;
        A7 : IN std_logic;
        A6 : IN std_logic;
        A5 : IN std_logic;
        A4 : IN std_logic;
        A3 : IN std_logic;
        A2 : IN std_logic;
        A1 : IN std_logic;
        A0 : IN std_logic;
        CO : OUT std_logic;
        Z7 : OUT std_logic;
        Z6 : OUT std_logic;
        Z5 : OUT std_logic;
        Z4 : OUT std_logic;
        Z3 : OUT std_logic;
        Z2 : OUT std_logic;
        Z1 : OUT std_logic;
        Z0 : OUT std_logic
    );
END ADDH8A;


ARCHITECTURE lattice_arch OF ADDH8A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, G012,
	 G345, P345 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => G012);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B4);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B5);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => A3);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N40, A1 => G012);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => B3, A1 => UQVN_N43);
UQVB_B7 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N3);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N37, A1 => B4, A2 => UQVN_N40);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N41, A1 => B3, A2 => G012);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => A3, A1 => UQVN_N41, A2 => G012);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B4, A1 => UQVN_N40, A2 => UQVN_N43);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N37, A1 => B4, A2 => UQVN_N43);
UQVB_B14 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N8);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A3, A1 => UQVN_N41, A2 => B3);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => A3, A1 => A4, A2 => A5, 
	A3 => B3);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A4, A1 => A5, A2 => B4);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => A3, A1 => A5, A2 => B3, 
	A3 => B4);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A5, A1 => B5);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => A3, A1 => A4, A2 => B3, 
	A3 => B5);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => A4, A1 => B4, A2 => B5);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => A3, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B24 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16, A6 => UQVN_N17);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N37, A1 => UQVN_N40);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N38, A1 => UQVN_N41);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N39, A1 => UQVN_N42);
UQVB_B28 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N20, A1 => UQVN_N18, A2 => UQVN_N19);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => B3);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A4);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A5);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N34);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N41, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N38, A1 => UQVN_N40, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N37, A1 => UQVN_N38, A2 => B5, 
	A3 => UQVN_N43);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => B3, A1 => B4, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => A3, A1 => B4, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A4, A1 => B3, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => A3, A1 => A4, A2 => UQVN_N42, 
	A3 => G012);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => A3, A1 => B3, A2 => B4, 
	A3 => UQVN_N42);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => A4, A1 => B4, A2 => UQVN_N42);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => A3, A1 => A4, A2 => B3, 
	A3 => UQVN_N42);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N37, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => B5);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N38, A1 => UQVN_N41, A2 => B5);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N37, A1 => UQVN_N38, A2 => UQVN_N40, 
	A3 => B5);
UQVB_B47 : OR12
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N28, A5 => UQVN_N27, A6 => UQVN_N26, 
	A7 => UQVN_N25, A8 => UQVN_N24, A9 => UQVN_N23, A10 => UQVN_N22, 
	A11 => UQVN_N21);
UQVB_B48 : OR3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N33, A1 => UQVN_N35, A2 => UQVN_N36);
UQVB_B49 : AND2
	PORT MAP (Z0 => UQVN_N44, A0 => P345, A1 => G012);
UQVB_B50 : OR2
	PORT MAP (Z0 => UQVN_N91, A0 => G345, A1 => UQVN_N44);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => B1);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => A0);
UQVB_B53 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B54 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N48);
UQVB_B55 : AND3
	PORT MAP (Z0 => UQVN_N47, A0 => A0, A1 => UQVN_N68, A2 => B0);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N52, A0 => A0, A1 => A1, A2 => A2, 
	A3 => B0);
UQVB_B57 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => A1, A1 => A2, A2 => B1);
UQVB_B58 : AND4
	PORT MAP (Z0 => UQVN_N50, A0 => A0, A1 => A2, A2 => B0, 
	A3 => B1);
UQVB_B59 : AND2
	PORT MAP (Z0 => UQVN_N49, A0 => A2, A1 => B2);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N53, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B2);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N54, A0 => A1, A1 => B1, A2 => B2);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N55, A0 => A0, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B63 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N52, A1 => UQVN_N51, A2 => UQVN_N50, 
	A3 => UQVN_N49, A4 => UQVN_N53, A5 => UQVN_N54, A6 => UQVN_N55);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => B0);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => A1);
UQVB_B66 : AND2
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N65, A1 => B1);
UQVB_B67 : AND2
	PORT MAP (Z0 => UQVN_N45, A0 => B1, A1 => UQVN_N67);
UQVB_B68 : OR3
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N46, A1 => UQVN_N45, A2 => UQVN_N47);
UQVB_B69 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => B2);
UQVB_B70 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N60);
UQVB_B71 : AND4
	PORT MAP (Z0 => UQVN_N59, A0 => A0, A1 => B0, A2 => B1, 
	A3 => UQVN_N69);
UQVB_B72 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => A1, A1 => B1, A2 => UQVN_N69);
UQVB_B73 : AND4
	PORT MAP (Z0 => UQVN_N57, A0 => A0, A1 => A1, A2 => B0, 
	A3 => UQVN_N69);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N66, A1 => UQVN_N68, A2 => B2);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N67, A1 => UQVN_N68, A2 => B2);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N65, A1 => UQVN_N68, A2 => B2);
UQVB_B77 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N66, A1 => UQVN_N67, A2 => B2);
UQVB_B78 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N65, A1 => UQVN_N66, A2 => B2);
UQVB_B79 : OR8
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N64, A1 => UQVN_N63, A2 => UQVN_N62, 
	A3 => UQVN_N61, A4 => UQVN_N59, A5 => UQVN_N58, A6 => UQVN_N57, 
	A7 => UQVN_N56);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N90, A0 => UQVN_N91);
UQVB_B81 : AND3
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N91, A1 => A7, A2 => A6);
UQVB_B82 : AND3
	PORT MAP (Z0 => UQVN_N71, A0 => UQVN_N91, A1 => A7, A2 => B6);
UQVB_B83 : AND3
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N91, A1 => A6, A2 => B7);
UQVB_B84 : AND3
	PORT MAP (Z0 => UQVN_N73, A0 => UQVN_N91, A1 => B7, A2 => B6);
UQVB_B85 : AND3
	PORT MAP (Z0 => UQVN_N74, A0 => A7, A1 => A6, A2 => B6);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N76, A0 => A6, A1 => B7, A2 => B6);
UQVB_B87 : AND2
	PORT MAP (Z0 => UQVN_N75, A0 => A7, A1 => B7);
UQVB_B88 : OR7
	PORT MAP (Z0 => CO, A0 => UQVN_N72, A1 => UQVN_N71, A2 => UQVN_N70, 
	A3 => UQVN_N73, A4 => UQVN_N74, A5 => UQVN_N76, A6 => UQVN_N75);
UQVB_B89 : AND3
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N87, A1 => B7, A2 => UQVN_N90);
UQVB_B90 : AND3
	PORT MAP (Z0 => UQVN_N78, A0 => B7, A1 => UQVN_N88, A2 => UQVN_N90);
UQVB_B91 : AND3
	PORT MAP (Z0 => UQVN_N79, A0 => A6, A1 => UQVN_N89, A2 => UQVN_N91);
UQVB_B92 : AND3
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N89, A1 => B6, A2 => UQVN_N91);
UQVB_B93 : AND3
	PORT MAP (Z0 => UQVN_N81, A0 => UQVN_N87, A1 => B7, A2 => UQVN_N88);
UQVB_B94 : AND3
	PORT MAP (Z0 => UQVN_N82, A0 => A6, A1 => UQVN_N89, A2 => B6);
UQVB_B95 : OR6
	PORT MAP (Z0 => UQVN_N83, A0 => UQVN_N77, A1 => UQVN_N78, A2 => UQVN_N79, 
	A3 => UQVN_N80, A4 => UQVN_N81, A5 => UQVN_N82);
UQVB_B96 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N83);
UQVB_B97 : INV
	PORT MAP (ZN0 => UQVN_N88, A0 => B6);
UQVB_B98 : INV
	PORT MAP (ZN0 => UQVN_N89, A0 => B7);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N87, A0 => A6);
UQVB_B100 : XOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N84);
UQVB_B101 : AND2
	PORT MAP (Z0 => UQVN_N85, A0 => UQVN_N91, A1 => UQVN_N88);
UQVB_B102 : OR2
	PORT MAP (Z0 => UQVN_N84, A0 => UQVN_N85, A1 => UQVN_N86);
UQVB_B103 : AND2
	PORT MAP (Z0 => UQVN_N86, A0 => UQVN_N90, A1 => B6);
END lattice_arch;
-- VHDL netlist for BI11
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI11 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BI11;


ARCHITECTURE lattice_arch OF BI11 IS

  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BI14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI14 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BI14;


ARCHITECTURE lattice_arch OF BI14 IS

  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => A2, OE => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BI18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI18 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BI18;


ARCHITECTURE lattice_arch OF BI18 IS

  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => A2, OE => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => A0, OE => OE);
UQVB_B5 : XBIDI1
	PORT MAP (Z0 => Z4, XB0 => XB4, A0 => A4, OE => OE);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => Z5, XB0 => XB5, A0 => A5, OE => OE);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z6, XB0 => XB6, A0 => A6, OE => OE);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => Z7, XB0 => XB7, A0 => A7, OE => OE);
END lattice_arch;
-- VHDL netlist for BI21
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI21 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BI21;


ARCHITECTURE lattice_arch OF BI21 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => UQVN_N1, OE => OE);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
END lattice_arch;
-- VHDL netlist for BI24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BI24;


ARCHITECTURE lattice_arch OF BI24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => UQVN_N1, OE => OE);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => UQVN_N2, OE => OE);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A2);
UQVB_B5 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => UQVN_N3, OE => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A1);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => UQVN_N4, OE => OE);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
END lattice_arch;
-- VHDL netlist for BI28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI28 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BI28;


ARCHITECTURE lattice_arch OF BI28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => UQVN_N1, OE => OE);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => UQVN_N2, OE => OE);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A2);
UQVB_B5 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => UQVN_N3, OE => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A1);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => UQVN_N4, OE => OE);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => Z4, XB0 => XB4, A0 => UQVN_N5, OE => OE);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A4);
UQVB_B11 : XBIDI1
	PORT MAP (Z0 => Z5, XB0 => XB5, A0 => UQVN_N6, OE => OE);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A5);
UQVB_B13 : XBIDI1
	PORT MAP (Z0 => Z6, XB0 => XB6, A0 => UQVN_N7, OE => OE);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A6);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => Z7, XB0 => XB7, A0 => UQVN_N8, OE => OE);
UQVB_B16 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A7);
END lattice_arch;
-- VHDL netlist for BI31
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI31 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BI31;


ARCHITECTURE lattice_arch OF BI31 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => A0, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
END lattice_arch;
-- VHDL netlist for BI34
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI34 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BI34;


ARCHITECTURE lattice_arch OF BI34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => A3, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => A2, OE => UQVN_N2);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B5 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => A1, OE => UQVN_N3);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => A0, OE => UQVN_N4);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
END lattice_arch;
-- VHDL netlist for BI38
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI38 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BI38;


ARCHITECTURE lattice_arch OF BI38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => A3, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => A2, OE => UQVN_N2);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B5 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => A1, OE => UQVN_N3);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => A0, OE => UQVN_N4);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => Z4, XB0 => XB4, A0 => A4, OE => UQVN_N5);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => OE);
UQVB_B11 : XBIDI1
	PORT MAP (Z0 => Z5, XB0 => XB5, A0 => A5, OE => UQVN_N6);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B13 : XBIDI1
	PORT MAP (Z0 => Z6, XB0 => XB6, A0 => A6, OE => UQVN_N7);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => OE);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => Z7, XB0 => XB7, A0 => A7, OE => UQVN_N8);
UQVB_B16 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
END lattice_arch;
-- VHDL netlist for BI41
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI41 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BI41;


ARCHITECTURE lattice_arch OF BI41 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => UQVN_N2, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A0);
END lattice_arch;
-- VHDL netlist for BI44
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BI44;


ARCHITECTURE lattice_arch OF BI44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => UQVN_N2, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A3);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => UQVN_N4, OE => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => UQVN_N6, OE => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => OE);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A1);
UQVB_B10 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => UQVN_N8, OE => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => OE);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A0);
END lattice_arch;
-- VHDL netlist for BI48
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BI48 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BI48;


ARCHITECTURE lattice_arch OF BI48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XBIDI1
	PORT MAP (Z0 => Z3, XB0 => XB3, A0 => UQVN_N2, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A3);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => Z2, XB0 => XB2, A0 => UQVN_N4, OE => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XBIDI1
	PORT MAP (Z0 => Z1, XB0 => XB1, A0 => UQVN_N6, OE => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => OE);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A1);
UQVB_B10 : XBIDI1
	PORT MAP (Z0 => Z0, XB0 => XB0, A0 => UQVN_N8, OE => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => OE);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A0);
UQVB_B13 : XBIDI1
	PORT MAP (Z0 => Z4, XB0 => XB4, A0 => UQVN_N10, OE => UQVN_N9);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A4);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => Z5, XB0 => XB5, A0 => UQVN_N12, OE => UQVN_N11);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => OE);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => A5);
UQVB_B19 : XBIDI1
	PORT MAP (Z0 => Z6, XB0 => XB6, A0 => UQVN_N14, OE => UQVN_N13);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => OE);
UQVB_B21 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => A6);
UQVB_B22 : XBIDI1
	PORT MAP (Z0 => Z7, XB0 => XB7, A0 => UQVN_N16, OE => UQVN_N15);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => OE);
UQVB_B24 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => A7);
END lattice_arch;
-- VHDL netlist for BIID11
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID11 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID11;


ARCHITECTURE lattice_arch OF BIID11 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID14 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID14;


ARCHITECTURE lattice_arch OF BIID14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B3 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB2, A0 => A2, OE => OE);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, CLK => CLK);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, CLK => CLK);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID18 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID18;


ARCHITECTURE lattice_arch OF BIID18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB7, A0 => A7, OE => OE);
UQVB_B3 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB6, A0 => A6, OE => OE);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N3, CLK => CLK);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB5, A0 => A5, OE => OE);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N4, CLK => CLK);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB4, A0 => A4, OE => OE);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N5, CLK => CLK);
UQVB_B10 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB0, A0 => A0, OE => OE);
UQVB_B11 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N6, CLK => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N7, CLK => CLK);
UQVB_B14 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B15 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N8, CLK => CLK);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB2, A0 => A2, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID21
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID21 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID21;


ARCHITECTURE lattice_arch OF BIID21 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => UQVN_N1, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID24;


ARCHITECTURE lattice_arch OF BIID24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => UQVN_N1, OE => OE);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N4, CLK => CLK);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A2);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB2, A0 => UQVN_N3, OE => OE);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N6, CLK => CLK);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A1);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB1, A0 => UQVN_N5, OE => OE);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N8, CLK => CLK);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A0);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB0, A0 => UQVN_N7, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID28 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID28;


ARCHITECTURE lattice_arch OF BIID28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => UQVN_N1, OE => OE);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N4, CLK => CLK);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A6);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB6, A0 => UQVN_N3, OE => OE);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N6, CLK => CLK);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A5);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB5, A0 => UQVN_N5, OE => OE);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N8, CLK => CLK);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A4);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB4, A0 => UQVN_N7, OE => OE);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N10, CLK => CLK);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => A0);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => UQVN_N10, XB0 => XB0, A0 => UQVN_N9, OE => OE);
UQVB_B16 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N12, CLK => CLK);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => A1);
UQVB_B18 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB1, A0 => UQVN_N11, OE => OE);
UQVB_B19 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N14, CLK => CLK);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A3);
UQVB_B21 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB3, A0 => UQVN_N13, OE => OE);
UQVB_B22 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N16, CLK => CLK);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => A2);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N16, XB0 => XB2, A0 => UQVN_N15, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID31
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID31 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID31;


ARCHITECTURE lattice_arch OF BIID31 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB0, A0 => A0, OE => UQVN_N2);
END lattice_arch;
-- VHDL netlist for BIID34
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID34 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID34;


ARCHITECTURE lattice_arch OF BIID34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB3, A0 => A3, OE => UQVN_N2);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N3, CLK => CLK);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB2, A0 => A2, OE => UQVN_N4);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N5, CLK => CLK);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB1, A0 => A1, OE => UQVN_N6);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N7, CLK => CLK);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB0, A0 => A0, OE => UQVN_N8);
END lattice_arch;
-- VHDL netlist for BIID38
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID38 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID38;


ARCHITECTURE lattice_arch OF BIID38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB7, A0 => A7, OE => UQVN_N2);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N3, CLK => CLK);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB6, A0 => A6, OE => UQVN_N4);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N5, CLK => CLK);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB5, A0 => A5, OE => UQVN_N6);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N7, CLK => CLK);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB4, A0 => A4, OE => UQVN_N8);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N9, CLK => CLK);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => OE);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => UQVN_N9, XB0 => XB0, A0 => A0, OE => UQVN_N10);
UQVB_B16 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N11, CLK => CLK);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B18 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB1, A0 => A1, OE => UQVN_N12);
UQVB_B19 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N13, CLK => CLK);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => OE);
UQVB_B21 : XBIDI1
	PORT MAP (Z0 => UQVN_N13, XB0 => XB3, A0 => A3, OE => UQVN_N14);
UQVB_B22 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N15, CLK => CLK);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => OE);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB2, A0 => A2, OE => UQVN_N16);
END lattice_arch;
-- VHDL netlist for BIID41
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID41 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID41;


ARCHITECTURE lattice_arch OF BIID41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => UQVN_N1, OE => UQVN_N3);
END lattice_arch;
-- VHDL netlist for BIID44
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID44;


ARCHITECTURE lattice_arch OF BIID44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => UQVN_N1, OE => UQVN_N3);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, CLK => CLK);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB2, A0 => UQVN_N4, OE => UQVN_N6);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N8, CLK => CLK);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A1);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB1, A0 => UQVN_N7, OE => UQVN_N9);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N11, CLK => CLK);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A0);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB0, A0 => UQVN_N10, OE => UQVN_N12);
END lattice_arch;
-- VHDL netlist for BIID48
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID48 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID48;


ARCHITECTURE lattice_arch OF BIID48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, CLK => CLK);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => UQVN_N1, OE => UQVN_N3);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N5, CLK => CLK);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB6, A0 => UQVN_N4, OE => UQVN_N6);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N8, CLK => CLK);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A5);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB5, A0 => UQVN_N7, OE => UQVN_N9);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N11, CLK => CLK);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A4);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB4, A0 => UQVN_N10, OE => UQVN_N12);
UQVB_B17 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B19 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => OE);
UQVB_B20 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB0, A0 => UQVN_N13, OE => UQVN_N15);
UQVB_B21 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N17, CLK => CLK);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => A1);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N18, A0 => OE);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N17, XB0 => XB1, A0 => UQVN_N16, OE => UQVN_N18);
UQVB_B25 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N20, CLK => CLK);
UQVB_B26 : XINV
	PORT MAP (ZN0 => UQVN_N19, A0 => A3);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N21, A0 => OE);
UQVB_B28 : XBIDI1
	PORT MAP (Z0 => UQVN_N20, XB0 => XB3, A0 => UQVN_N19, OE => UQVN_N21);
UQVB_B29 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N23, CLK => CLK);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => A2);
UQVB_B31 : XINV
	PORT MAP (ZN0 => UQVN_N24, A0 => OE);
UQVB_B32 : XBIDI1
	PORT MAP (Z0 => UQVN_N23, XB0 => XB2, A0 => UQVN_N22, OE => UQVN_N24);
END lattice_arch;
-- VHDL netlist for BIID51
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID51 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID51;


ARCHITECTURE lattice_arch OF BIID51 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => CLK);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID54
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID54 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID54;


ARCHITECTURE lattice_arch OF BIID54 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => CLK);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N4, CLK => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => CLK);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB2, A0 => A2, OE => OE);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N6, CLK => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => CLK);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N8, CLK => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID58
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID58 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID58;


ARCHITECTURE lattice_arch OF BIID58 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, CLK => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => CLK);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => A7, OE => OE);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N4, CLK => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => CLK);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB6, A0 => A6, OE => OE);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N6, CLK => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => CLK);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB5, A0 => A5, OE => OE);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N8, CLK => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB4, A0 => A4, OE => OE);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N10, CLK => UQVN_N9);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => CLK);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => UQVN_N10, XB0 => XB0, A0 => A0, OE => OE);
UQVB_B16 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N12, CLK => UQVN_N11);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => CLK);
UQVB_B18 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B19 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N14, CLK => UQVN_N13);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => CLK);
UQVB_B21 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B22 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N16, CLK => UQVN_N15);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => CLK);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N16, XB0 => XB2, A0 => A2, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID61
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID61 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID61;


ARCHITECTURE lattice_arch OF BIID61 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N3, CLK => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB0, A0 => UQVN_N1, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID64
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID64 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID64;


ARCHITECTURE lattice_arch OF BIID64 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, CLK => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB3, A0 => UQVN_N1, OE => OE);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => UQVN_N5);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => CLK);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB2, A0 => UQVN_N4, OE => OE);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N9, CLK => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A1);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N9, XB0 => XB1, A0 => UQVN_N7, OE => OE);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N12, CLK => UQVN_N11);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A0);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => CLK);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB0, A0 => UQVN_N10, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID68
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID68 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID68;


ARCHITECTURE lattice_arch OF BIID68 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N3, CLK => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB7, A0 => UQVN_N1, OE => OE);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N6, CLK => UQVN_N5);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => CLK);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB6, A0 => UQVN_N4, OE => OE);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N9, CLK => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A5);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N9, XB0 => XB5, A0 => UQVN_N7, OE => OE);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N12, CLK => UQVN_N11);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A4);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => CLK);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB4, A0 => UQVN_N10, OE => OE);
UQVB_B17 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N15, CLK => UQVN_N14);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B19 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => CLK);
UQVB_B20 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB0, A0 => UQVN_N13, OE => OE);
UQVB_B21 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N18, CLK => UQVN_N17);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => A1);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N17, A0 => CLK);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N18, XB0 => XB1, A0 => UQVN_N16, OE => OE);
UQVB_B25 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N21, CLK => UQVN_N20);
UQVB_B26 : XINV
	PORT MAP (ZN0 => UQVN_N19, A0 => A3);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N20, A0 => CLK);
UQVB_B28 : XBIDI1
	PORT MAP (Z0 => UQVN_N21, XB0 => XB3, A0 => UQVN_N19, OE => OE);
UQVB_B29 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N24, CLK => UQVN_N23);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => A2);
UQVB_B31 : XINV
	PORT MAP (ZN0 => UQVN_N23, A0 => CLK);
UQVB_B32 : XBIDI1
	PORT MAP (Z0 => UQVN_N24, XB0 => XB2, A0 => UQVN_N22, OE => OE);
END lattice_arch;
-- VHDL netlist for BIID71
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID71 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID71;


ARCHITECTURE lattice_arch OF BIID71 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => A0, OE => UQVN_N3);
END lattice_arch;
-- VHDL netlist for BIID74
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID74 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID74;


ARCHITECTURE lattice_arch OF BIID74 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => A3, OE => UQVN_N3);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, CLK => UQVN_N4);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => CLK);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB2, A0 => A2, OE => UQVN_N6);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N8, CLK => UQVN_N7);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB1, A0 => A1, OE => UQVN_N9);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N11, CLK => UQVN_N10);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => CLK);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB0, A0 => A0, OE => UQVN_N12);
END lattice_arch;
-- VHDL netlist for BIID78
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID78 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID78;


ARCHITECTURE lattice_arch OF BIID78 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, CLK => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => A7, OE => UQVN_N3);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N5, CLK => UQVN_N4);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => CLK);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB6, A0 => A6, OE => UQVN_N6);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N8, CLK => UQVN_N7);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => CLK);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB5, A0 => A5, OE => UQVN_N9);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N11, CLK => UQVN_N10);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => CLK);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB4, A0 => A4, OE => UQVN_N12);
UQVB_B17 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => UQVN_N13);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => OE);
UQVB_B19 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => CLK);
UQVB_B20 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB0, A0 => A0, OE => UQVN_N15);
UQVB_B21 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N17, CLK => UQVN_N16);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N18, A0 => OE);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => CLK);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N17, XB0 => XB1, A0 => A1, OE => UQVN_N18);
UQVB_B25 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N20, CLK => UQVN_N19);
UQVB_B26 : XINV
	PORT MAP (ZN0 => UQVN_N21, A0 => OE);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N19, A0 => CLK);
UQVB_B28 : XBIDI1
	PORT MAP (Z0 => UQVN_N20, XB0 => XB3, A0 => A3, OE => UQVN_N21);
UQVB_B29 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N23, CLK => UQVN_N22);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N24, A0 => OE);
UQVB_B31 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => CLK);
UQVB_B32 : XBIDI1
	PORT MAP (Z0 => UQVN_N23, XB0 => XB2, A0 => A2, OE => UQVN_N24);
END lattice_arch;
-- VHDL netlist for BIID81
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID81 IS 
    PORT (
        A0 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIID81;


ARCHITECTURE lattice_arch OF BIID81 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N3, CLK => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB0, A0 => UQVN_N1, OE => UQVN_N4);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
END lattice_arch;
-- VHDL netlist for BIID84
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID84 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIID84;


ARCHITECTURE lattice_arch OF BIID84 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, CLK => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB3, A0 => UQVN_N1, OE => UQVN_N4);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N7, CLK => UQVN_N6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A2);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => CLK);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB2, A0 => UQVN_N5, OE => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B11 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N11, CLK => UQVN_N10);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => A1);
UQVB_B13 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => CLK);
UQVB_B14 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB1, A0 => UQVN_N9, OE => UQVN_N12);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N15, CLK => UQVN_N14);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => CLK);
UQVB_B19 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB0, A0 => UQVN_N13, OE => UQVN_N16);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => OE);
END lattice_arch;
-- VHDL netlist for BIID88
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIID88 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        CLK : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIID88;


ARCHITECTURE lattice_arch OF BIID88 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N3, CLK => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB7, A0 => UQVN_N1, OE => UQVN_N4);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N7, CLK => UQVN_N6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A6);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => CLK);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB6, A0 => UQVN_N5, OE => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B11 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N11, CLK => UQVN_N10);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => A5);
UQVB_B13 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => CLK);
UQVB_B14 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB5, A0 => UQVN_N9, OE => UQVN_N12);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N15, CLK => UQVN_N14);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A4);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => CLK);
UQVB_B19 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB4, A0 => UQVN_N13, OE => UQVN_N16);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => OE);
UQVB_B21 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N19, CLK => UQVN_N18);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N17, A0 => A0);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N18, A0 => CLK);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N19, XB0 => XB0, A0 => UQVN_N17, OE => UQVN_N20);
UQVB_B25 : XINV
	PORT MAP (ZN0 => UQVN_N20, A0 => OE);
UQVB_B26 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N23, CLK => UQVN_N22);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N21, A0 => A1);
UQVB_B28 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => CLK);
UQVB_B29 : XBIDI1
	PORT MAP (Z0 => UQVN_N23, XB0 => XB1, A0 => UQVN_N21, OE => UQVN_N24);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N24, A0 => OE);
UQVB_B31 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N27, CLK => UQVN_N26);
UQVB_B32 : XINV
	PORT MAP (ZN0 => UQVN_N25, A0 => A3);
UQVB_B33 : XINV
	PORT MAP (ZN0 => UQVN_N26, A0 => CLK);
UQVB_B34 : XBIDI1
	PORT MAP (Z0 => UQVN_N27, XB0 => XB3, A0 => UQVN_N25, OE => UQVN_N28);
UQVB_B35 : XINV
	PORT MAP (ZN0 => UQVN_N28, A0 => OE);
UQVB_B36 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N31, CLK => UQVN_N30);
UQVB_B37 : XINV
	PORT MAP (ZN0 => UQVN_N29, A0 => A2);
UQVB_B38 : XINV
	PORT MAP (ZN0 => UQVN_N30, A0 => CLK);
UQVB_B39 : XBIDI1
	PORT MAP (Z0 => UQVN_N31, XB0 => XB2, A0 => UQVN_N29, OE => UQVN_N32);
UQVB_B40 : XINV
	PORT MAP (ZN0 => UQVN_N32, A0 => OE);
END lattice_arch;
-- VHDL netlist for BIIL11
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL11 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL11;


ARCHITECTURE lattice_arch OF BIIL11 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, G => G);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL14 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL14;


ARCHITECTURE lattice_arch OF BIIL14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, G => G);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B3 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, G => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB2, A0 => A2, OE => OE);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, G => G);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, G => G);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL18 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL18;


ARCHITECTURE lattice_arch OF BIIL18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N1, G => G);
UQVB_B2 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB7, A0 => A7, OE => OE);
UQVB_B3 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N2, G => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB6, A0 => A6, OE => OE);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N3, G => G);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB5, A0 => A5, OE => OE);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N4, G => G);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB4, A0 => A4, OE => OE);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N5, G => G);
UQVB_B10 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB0, A0 => A0, OE => OE);
UQVB_B11 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N6, G => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N7, G => G);
UQVB_B14 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B15 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N8, G => G);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB2, A0 => A2, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL21
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL21 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL21;


ARCHITECTURE lattice_arch OF BIIL21 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => UQVN_N1, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL24;


ARCHITECTURE lattice_arch OF BIIL24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => UQVN_N1, OE => OE);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N4, G => G);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A2);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB2, A0 => UQVN_N3, OE => OE);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N6, G => G);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A1);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB1, A0 => UQVN_N5, OE => OE);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N8, G => G);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A0);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB0, A0 => UQVN_N7, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL28 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL28;


ARCHITECTURE lattice_arch OF BIIL28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => UQVN_N1, OE => OE);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N4, G => G);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A6);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB6, A0 => UQVN_N3, OE => OE);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N6, G => G);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A5);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB5, A0 => UQVN_N5, OE => OE);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N8, G => G);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A4);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB4, A0 => UQVN_N7, OE => OE);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N10, G => G);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => A0);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => UQVN_N10, XB0 => XB0, A0 => UQVN_N9, OE => OE);
UQVB_B16 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N12, G => G);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => A1);
UQVB_B18 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB1, A0 => UQVN_N11, OE => OE);
UQVB_B19 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N14, G => G);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A3);
UQVB_B21 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB3, A0 => UQVN_N13, OE => OE);
UQVB_B22 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N16, G => G);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => A2);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N16, XB0 => XB2, A0 => UQVN_N15, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL31
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL31 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL31;


ARCHITECTURE lattice_arch OF BIIL31 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB0, A0 => A0, OE => UQVN_N2);
END lattice_arch;
-- VHDL netlist for BIIL34
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL34 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL34;


ARCHITECTURE lattice_arch OF BIIL34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB3, A0 => A3, OE => UQVN_N2);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N3, G => G);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB2, A0 => A2, OE => UQVN_N4);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N5, G => G);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB1, A0 => A1, OE => UQVN_N6);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N7, G => G);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB0, A0 => A0, OE => UQVN_N8);
END lattice_arch;
-- VHDL netlist for BIIL38
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL38 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL38;


ARCHITECTURE lattice_arch OF BIIL38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N1, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N1, XB0 => XB7, A0 => A7, OE => UQVN_N2);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N3, G => G);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB6, A0 => A6, OE => UQVN_N4);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N5, G => G);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB5, A0 => A5, OE => UQVN_N6);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N7, G => G);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB4, A0 => A4, OE => UQVN_N8);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N9, G => G);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => OE);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => UQVN_N9, XB0 => XB0, A0 => A0, OE => UQVN_N10);
UQVB_B16 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N11, G => G);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B18 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB1, A0 => A1, OE => UQVN_N12);
UQVB_B19 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N13, G => G);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => OE);
UQVB_B21 : XBIDI1
	PORT MAP (Z0 => UQVN_N13, XB0 => XB3, A0 => A3, OE => UQVN_N14);
UQVB_B22 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N15, G => G);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => OE);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB2, A0 => A2, OE => UQVN_N16);
END lattice_arch;
-- VHDL netlist for BIIL41
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL41 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL41;


ARCHITECTURE lattice_arch OF BIIL41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => UQVN_N1, OE => UQVN_N3);
END lattice_arch;
-- VHDL netlist for BIIL44
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL44;


ARCHITECTURE lattice_arch OF BIIL44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => UQVN_N1, OE => UQVN_N3);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, G => G);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB2, A0 => UQVN_N4, OE => UQVN_N6);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N8, G => G);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A1);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB1, A0 => UQVN_N7, OE => UQVN_N9);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N11, G => G);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A0);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB0, A0 => UQVN_N10, OE => UQVN_N12);
END lattice_arch;
-- VHDL netlist for BIIL48
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL48 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL48;


ARCHITECTURE lattice_arch OF BIIL48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, G => G);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => UQVN_N1, OE => UQVN_N3);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N5, G => G);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB6, A0 => UQVN_N4, OE => UQVN_N6);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N8, G => G);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A5);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB5, A0 => UQVN_N7, OE => UQVN_N9);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N11, G => G);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A4);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB4, A0 => UQVN_N10, OE => UQVN_N12);
UQVB_B17 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, G => G);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B19 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => OE);
UQVB_B20 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB0, A0 => UQVN_N13, OE => UQVN_N15);
UQVB_B21 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N17, G => G);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => A1);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N18, A0 => OE);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N17, XB0 => XB1, A0 => UQVN_N16, OE => UQVN_N18);
UQVB_B25 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N20, G => G);
UQVB_B26 : XINV
	PORT MAP (ZN0 => UQVN_N19, A0 => A3);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N21, A0 => OE);
UQVB_B28 : XBIDI1
	PORT MAP (Z0 => UQVN_N20, XB0 => XB3, A0 => UQVN_N19, OE => UQVN_N21);
UQVB_B29 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N23, G => G);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => A2);
UQVB_B31 : XINV
	PORT MAP (ZN0 => UQVN_N24, A0 => OE);
UQVB_B32 : XBIDI1
	PORT MAP (Z0 => UQVN_N23, XB0 => XB2, A0 => UQVN_N22, OE => UQVN_N24);
END lattice_arch;
-- VHDL netlist for BIIL51
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL51 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL51;


ARCHITECTURE lattice_arch OF BIIL51 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, G => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => G);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL54
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL54 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL54;


ARCHITECTURE lattice_arch OF BIIL54 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, G => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => G);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N4, G => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => G);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB2, A0 => A2, OE => OE);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N6, G => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N8, G => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL58
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL58 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL58;


ARCHITECTURE lattice_arch OF BIIL58 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, G => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => G);
UQVB_B3 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => A7, OE => OE);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N4, G => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => G);
UQVB_B6 : XBIDI1
	PORT MAP (Z0 => UQVN_N4, XB0 => XB6, A0 => A6, OE => OE);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N6, G => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB5, A0 => A5, OE => OE);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N8, G => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB4, A0 => A4, OE => OE);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N10, G => UQVN_N9);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => G);
UQVB_B15 : XBIDI1
	PORT MAP (Z0 => UQVN_N10, XB0 => XB0, A0 => A0, OE => OE);
UQVB_B16 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N12, G => UQVN_N11);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B18 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB1, A0 => A1, OE => OE);
UQVB_B19 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N14, G => UQVN_N13);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => G);
UQVB_B21 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB3, A0 => A3, OE => OE);
UQVB_B22 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N16, G => UQVN_N15);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => G);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N16, XB0 => XB2, A0 => A2, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL61
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL61 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL61;


ARCHITECTURE lattice_arch OF BIIL61 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N3, G => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB0, A0 => UQVN_N1, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL64
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL64 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL64;


ARCHITECTURE lattice_arch OF BIIL64 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, G => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB3, A0 => UQVN_N1, OE => OE);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, G => UQVN_N5);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB2, A0 => UQVN_N4, OE => OE);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N9, G => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A1);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N9, XB0 => XB1, A0 => UQVN_N7, OE => OE);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N12, G => UQVN_N11);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A0);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB0, A0 => UQVN_N10, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL68
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL68 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL68;


ARCHITECTURE lattice_arch OF BIIL68 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N3, G => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB7, A0 => UQVN_N1, OE => OE);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N6, G => UQVN_N5);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N6, XB0 => XB6, A0 => UQVN_N4, OE => OE);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N9, G => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A5);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N9, XB0 => XB5, A0 => UQVN_N7, OE => OE);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N12, G => UQVN_N11);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A4);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N12, XB0 => XB4, A0 => UQVN_N10, OE => OE);
UQVB_B17 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N15, G => UQVN_N14);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B19 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B20 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB0, A0 => UQVN_N13, OE => OE);
UQVB_B21 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N18, G => UQVN_N17);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => A1);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N17, A0 => G);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N18, XB0 => XB1, A0 => UQVN_N16, OE => OE);
UQVB_B25 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N21, G => UQVN_N20);
UQVB_B26 : XINV
	PORT MAP (ZN0 => UQVN_N19, A0 => A3);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N20, A0 => G);
UQVB_B28 : XBIDI1
	PORT MAP (Z0 => UQVN_N21, XB0 => XB3, A0 => UQVN_N19, OE => OE);
UQVB_B29 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N24, G => UQVN_N23);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => A2);
UQVB_B31 : XINV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B32 : XBIDI1
	PORT MAP (Z0 => UQVN_N24, XB0 => XB2, A0 => UQVN_N22, OE => OE);
END lattice_arch;
-- VHDL netlist for BIIL71
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL71 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL71;


ARCHITECTURE lattice_arch OF BIIL71 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, G => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB0, A0 => A0, OE => UQVN_N3);
END lattice_arch;
-- VHDL netlist for BIIL74
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL74 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL74;


ARCHITECTURE lattice_arch OF BIIL74 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, G => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB3, A0 => A3, OE => UQVN_N3);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, G => UQVN_N4);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB2, A0 => A2, OE => UQVN_N6);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N8, G => UQVN_N7);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB1, A0 => A1, OE => UQVN_N9);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N11, G => UQVN_N10);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => G);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB0, A0 => A0, OE => UQVN_N12);
END lattice_arch;
-- VHDL netlist for BIIL78
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL78 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL78;


ARCHITECTURE lattice_arch OF BIIL78 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, G => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N2, XB0 => XB7, A0 => A7, OE => UQVN_N3);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N5, G => UQVN_N4);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B8 : XBIDI1
	PORT MAP (Z0 => UQVN_N5, XB0 => XB6, A0 => A6, OE => UQVN_N6);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N8, G => UQVN_N7);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B12 : XBIDI1
	PORT MAP (Z0 => UQVN_N8, XB0 => XB5, A0 => A5, OE => UQVN_N9);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N11, G => UQVN_N10);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => G);
UQVB_B16 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB4, A0 => A4, OE => UQVN_N12);
UQVB_B17 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, G => UQVN_N13);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => OE);
UQVB_B19 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => G);
UQVB_B20 : XBIDI1
	PORT MAP (Z0 => UQVN_N14, XB0 => XB0, A0 => A0, OE => UQVN_N15);
UQVB_B21 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N17, G => UQVN_N16);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N18, A0 => OE);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => G);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N17, XB0 => XB1, A0 => A1, OE => UQVN_N18);
UQVB_B25 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N20, G => UQVN_N19);
UQVB_B26 : XINV
	PORT MAP (ZN0 => UQVN_N21, A0 => OE);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N19, A0 => G);
UQVB_B28 : XBIDI1
	PORT MAP (Z0 => UQVN_N20, XB0 => XB3, A0 => A3, OE => UQVN_N21);
UQVB_B29 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N23, G => UQVN_N22);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N24, A0 => OE);
UQVB_B31 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => G);
UQVB_B32 : XBIDI1
	PORT MAP (Z0 => UQVN_N23, XB0 => XB2, A0 => A2, OE => UQVN_N24);
END lattice_arch;
-- VHDL netlist for BIIL81
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL81 IS 
    PORT (
        A0 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
END BIIL81;


ARCHITECTURE lattice_arch OF BIIL81 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N3, G => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB0, A0 => UQVN_N1, OE => UQVN_N4);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
END lattice_arch;
-- VHDL netlist for BIIL84
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL84 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic
    );
END BIIL84;


ARCHITECTURE lattice_arch OF BIIL84 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, G => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB3, A0 => UQVN_N1, OE => UQVN_N4);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N7, G => UQVN_N6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A2);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB2, A0 => UQVN_N5, OE => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B11 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N11, G => UQVN_N10);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => A1);
UQVB_B13 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => G);
UQVB_B14 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB1, A0 => UQVN_N9, OE => UQVN_N12);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N15, G => UQVN_N14);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B19 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB0, A0 => UQVN_N13, OE => UQVN_N16);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => OE);
END lattice_arch;
-- VHDL netlist for BIIL88
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIIL88 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        G : IN std_logic;
        OE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        XB0 : INOUT std_logic;
        XB1 : INOUT std_logic;
        XB2 : INOUT std_logic;
        XB3 : INOUT std_logic;
        XB4 : INOUT std_logic;
        XB5 : INOUT std_logic;
        XB6 : INOUT std_logic;
        XB7 : INOUT std_logic
    );
END BIIL88;


ARCHITECTURE lattice_arch OF BIIL88 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


  COMPONENT XBIDI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        Z0 : OUT std_logic;
        XB0 : INOUT std_logic
    );
  END COMPONENT;

for all: XBIDI1 use  entity  lat_vhd.XBIDI1(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N3, G => UQVN_N2);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A7);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XBIDI1
	PORT MAP (Z0 => UQVN_N3, XB0 => XB7, A0 => UQVN_N1, OE => UQVN_N4);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B6 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N7, G => UQVN_N6);
UQVB_B7 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A6);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B9 : XBIDI1
	PORT MAP (Z0 => UQVN_N7, XB0 => XB6, A0 => UQVN_N5, OE => UQVN_N8);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
UQVB_B11 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N11, G => UQVN_N10);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => A5);
UQVB_B13 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => G);
UQVB_B14 : XBIDI1
	PORT MAP (Z0 => UQVN_N11, XB0 => XB5, A0 => UQVN_N9, OE => UQVN_N12);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => OE);
UQVB_B16 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N15, G => UQVN_N14);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => A4);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B19 : XBIDI1
	PORT MAP (Z0 => UQVN_N15, XB0 => XB4, A0 => UQVN_N13, OE => UQVN_N16);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => OE);
UQVB_B21 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N19, G => UQVN_N18);
UQVB_B22 : XINV
	PORT MAP (ZN0 => UQVN_N17, A0 => A0);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N18, A0 => G);
UQVB_B24 : XBIDI1
	PORT MAP (Z0 => UQVN_N19, XB0 => XB0, A0 => UQVN_N17, OE => UQVN_N20);
UQVB_B25 : XINV
	PORT MAP (ZN0 => UQVN_N20, A0 => OE);
UQVB_B26 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N23, G => UQVN_N22);
UQVB_B27 : XINV
	PORT MAP (ZN0 => UQVN_N21, A0 => A1);
UQVB_B28 : XINV
	PORT MAP (ZN0 => UQVN_N22, A0 => G);
UQVB_B29 : XBIDI1
	PORT MAP (Z0 => UQVN_N23, XB0 => XB1, A0 => UQVN_N21, OE => UQVN_N24);
UQVB_B30 : XINV
	PORT MAP (ZN0 => UQVN_N24, A0 => OE);
UQVB_B31 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N27, G => UQVN_N26);
UQVB_B32 : XINV
	PORT MAP (ZN0 => UQVN_N25, A0 => A3);
UQVB_B33 : XINV
	PORT MAP (ZN0 => UQVN_N26, A0 => G);
UQVB_B34 : XBIDI1
	PORT MAP (Z0 => UQVN_N27, XB0 => XB3, A0 => UQVN_N25, OE => UQVN_N28);
UQVB_B35 : XINV
	PORT MAP (ZN0 => UQVN_N28, A0 => OE);
UQVB_B36 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N31, G => UQVN_N30);
UQVB_B37 : XINV
	PORT MAP (ZN0 => UQVN_N29, A0 => A2);
UQVB_B38 : XINV
	PORT MAP (ZN0 => UQVN_N30, A0 => G);
UQVB_B39 : XBIDI1
	PORT MAP (Z0 => UQVN_N31, XB0 => XB2, A0 => UQVN_N29, OE => UQVN_N32);
UQVB_B40 : XINV
	PORT MAP (ZN0 => UQVN_N32, A0 => OE);
END lattice_arch;
-- VHDL netlist for BIN27
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY BIN27 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        EN : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic
    );
END BIN27;


ARCHITECTURE lattice_arch OF BIN27 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => A0);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => A1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => A2);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => EN, A1 => A1, A2 => UQVN_N35);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A3);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => EN, A1 => A3, A2 => UQVN_N37);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => EN, A1 => UQVN_N38, A2 => A2, 
	A3 => A0);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => EN, A1 => A2, A2 => A1);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => EN, A1 => UQVN_N38, A2 => A1);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => A3, A2 => UQVN_N37, 
	A3 => UQVN_N36);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35);
UQVB_B12 : OR6
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N4, A4 => UQVN_N5, A5 => UQVN_N6);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => EN, A1 => UQVN_N38, A2 => UQVN_N37);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => EN, A1 => UQVN_N38, A2 => A1, 
	A3 => A0);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => EN, A1 => A3, A2 => UQVN_N36, 
	A3 => A0);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => EN, A1 => UQVN_N38, A2 => UQVN_N36, 
	A3 => UQVN_N35);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => EN, A1 => A3, A2 => UQVN_N37, 
	A3 => UQVN_N35);
UQVB_B18 : OR5
	PORT MAP (Z0 => Z1, A0 => UQVN_N9, A1 => UQVN_N8, A2 => UQVN_N7, 
	A3 => UQVN_N10, A4 => UQVN_N11);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => EN, A1 => UQVN_N36, A2 => A0);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => EN, A1 => UQVN_N38, A2 => A2);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => EN, A1 => UQVN_N38, A2 => A0);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => EN, A1 => UQVN_N38, A2 => UQVN_N36);
UQVB_B23 : OR5
	PORT MAP (Z0 => Z2, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N15, A4 => UQVN_N16);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => EN, A1 => A3, A2 => UQVN_N36);
UQVB_B25 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => EN, A1 => A2, A2 => UQVN_N36, 
	A3 => A0);
UQVB_B26 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => EN, A1 => A2, A2 => A1, 
	A3 => UQVN_N35);
UQVB_B27 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => EN, A1 => UQVN_N37, A2 => A1, 
	A3 => A0);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => EN, A1 => UQVN_N38, A2 => UQVN_N37, 
	A3 => UQVN_N35);
UQVB_B29 : OR5
	PORT MAP (Z0 => Z3, A0 => UQVN_N19, A1 => UQVN_N18, A2 => UQVN_N17, 
	A3 => UQVN_N20, A4 => UQVN_N21);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => EN, A1 => A1, A2 => UQVN_N35);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => EN, A1 => A3, A2 => A2);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => EN, A1 => A3, A2 => A1);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35);
UQVB_B34 : OR4
	PORT MAP (Z0 => Z4, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N22, 
	A3 => UQVN_N25);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => EN, A1 => A3, A2 => UQVN_N37);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => EN, A1 => A3, A2 => A1);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => EN, A1 => UQVN_N38, A2 => A2, 
	A3 => UQVN_N36);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => EN, A1 => A2, A2 => A1, 
	A3 => UQVN_N35);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35);
UQVB_B40 : OR5
	PORT MAP (Z0 => Z5, A0 => UQVN_N28, A1 => UQVN_N27, A2 => UQVN_N26, 
	A3 => UQVN_N29, A4 => UQVN_N30);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => EN, A1 => A1, A2 => UQVN_N35);
UQVB_B42 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => EN, A1 => A3);
UQVB_B43 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => EN, A1 => A2, A2 => UQVN_N36);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => EN, A1 => UQVN_N37, A2 => A1, 
	A3 => A0);
UQVB_B45 : OR4
	PORT MAP (Z0 => Z6, A0 => UQVN_N33, A1 => UQVN_N32, A2 => UQVN_N31, 
	A3 => UQVN_N34);
END lattice_arch;
-- VHDL netlist for CBD11
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD11 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD11;


ARCHITECTURE lattice_arch OF CBD11 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => UQVN_N1);
UQVB_B3 : AND2
	PORT MAP (Z0 => CAO, A0 => UQVN_N2, A1 => CAI);
UQVB_B4 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N1);
UQVB_B5 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => CAI);
END lattice_arch;
-- VHDL netlist for CBD12
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD12 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD12;


ARCHITECTURE lattice_arch OF CBD12 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, QI0,
	 QI1, UQVN_N4, UQVN_N5 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => QI1);
UQVB_B5 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N4, A1 => UQVN_N5, A2 => CAI);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N4, A1 => CAI);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B9 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI);
UQVB_B10 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for CBD14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD14 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD14;


ARCHITECTURE lattice_arch OF CBD14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, QI0,
	 QI1, QI2, QI3, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => QI1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => QI2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => QI3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => CAI);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N9, A2 => CAI);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => CAI);
UQVB_B10 : AND5
	PORT MAP (Z0 => CAO, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => CAI);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B15 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B16 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => CAI);
UQVB_B18 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => QI1, A1 => UQVN_N1);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => UQVN_N6, A0 => QI2, A1 => UQVN_N2);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for CBD18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD18 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD18;


ARCHITECTURE lattice_arch OF CBD18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, QI0,
	 QI1, QI2, QI3, QI4,
	 QI5, QI6, QI7, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => QI1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => QI2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => QI3);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => QI4);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => QI5);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => QI6);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI7);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N16, A1 => CAI);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N16, A1 => UQVN_N17, A2 => CAI);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N16, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => CAI);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N16, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => CAI);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N16, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => CAI);
UQVB_B16 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N16, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => UQVN_N21, A6 => CAI);
UQVB_B17 : AND8
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N16, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => UQVN_N21, A6 => UQVN_N22, 
	A7 => CAI);
UQVB_B18 : AND9
	PORT MAP (Z0 => CAO, A0 => UQVN_N16, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => UQVN_N21, A6 => UQVN_N22, 
	A7 => UQVN_N23, A8 => CAI);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B27 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => QI0, A1 => CAI);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI1, A1 => UQVN_N1);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI2, A1 => UQVN_N2);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => QI3, A1 => UQVN_N3);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => QI4, A1 => UQVN_N4);
UQVB_B34 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => QI5, A1 => UQVN_N5);
UQVB_B36 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B37 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B38 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => QI6, A1 => UQVN_N6);
UQVB_B39 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => QI7, A1 => UQVN_N7);
UQVB_B40 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N15, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CBD21
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD21 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD21;


ARCHITECTURE lattice_arch OF CBD21 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => UQVN_N1);
UQVB_B3 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N4, A1 => CAI, A2 => EN);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => CAI, A1 => EN);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N1);
UQVB_B6 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => UQVN_N2);
END lattice_arch;
-- VHDL netlist for CBD22
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD22 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD22;


ARCHITECTURE lattice_arch OF CBD22 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 QI0, QI1, UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => QI1);
UQVB_B5 : AND4
	PORT MAP (Z0 => CAO, A0 => UQVN_N5, A1 => UQVN_N6, A2 => CAI, 
	A3 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => CAI, A2 => EN);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B10 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI0, A1 => UQVN_N1);
UQVB_B11 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI1, A1 => UQVN_N2);
END lattice_arch;
-- VHDL netlist for CBD24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD24 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD24;


ARCHITECTURE lattice_arch OF CBD24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 QI0, QI1, QI2, QI3,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => QI1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => QI2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => QI3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N9, A1 => CAI, A2 => EN);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N9, A1 => UQVN_N10, A2 => CAI, 
	A3 => EN);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N9, A1 => UQVN_N10, A2 => UQVN_N11, 
	A3 => CAI, A4 => EN);
UQVB_B11 : AND6
	PORT MAP (Z0 => CAO, A0 => UQVN_N9, A1 => UQVN_N10, A2 => UQVN_N11, 
	A3 => UQVN_N12, A4 => CAI, A5 => EN);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B16 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B17 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B18 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => UQVN_N1);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => UQVN_N6, A0 => QI1, A1 => UQVN_N2);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => QI2, A1 => UQVN_N3);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => UQVN_N4);
END lattice_arch;
-- VHDL netlist for CBD28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD28 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD28;


ARCHITECTURE lattice_arch OF CBD28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 QI0, QI1, QI2, QI3,
	 QI4, QI5, QI6, QI7,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => QI1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => QI2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => QI3);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => QI4);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => QI5);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI6);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI7);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N17, A1 => CAI, A2 => EN);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N17, A1 => UQVN_N18, A2 => CAI, 
	A3 => EN);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => UQVN_N18, A2 => UQVN_N19, 
	A3 => CAI, A4 => EN);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N17, A1 => UQVN_N18, A2 => UQVN_N19, 
	A3 => UQVN_N20, A4 => CAI, A5 => EN);
UQVB_B16 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N17, A1 => UQVN_N18, A2 => UQVN_N19, 
	A3 => UQVN_N20, A4 => UQVN_N21, A5 => CAI, A6 => EN);
UQVB_B17 : AND8
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N17, A1 => UQVN_N18, A2 => UQVN_N19, 
	A3 => UQVN_N20, A4 => UQVN_N21, A5 => UQVN_N22, A6 => CAI, 
	A7 => EN);
UQVB_B18 : AND9
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N17, A1 => UQVN_N18, A2 => UQVN_N19, 
	A3 => UQVN_N20, A4 => UQVN_N21, A5 => UQVN_N22, A6 => UQVN_N23, 
	A7 => CAI, A8 => EN);
UQVB_B19 : AND10
	PORT MAP (Z0 => CAO, A0 => UQVN_N17, A1 => UQVN_N18, A2 => UQVN_N19, 
	A3 => UQVN_N20, A4 => UQVN_N21, A5 => UQVN_N22, A6 => UQVN_N23, 
	A7 => UQVN_N24, A8 => CAI, A9 => EN);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI0, A1 => UQVN_N1);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI1, A1 => UQVN_N2);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => QI2, A1 => UQVN_N3);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => QI3, A1 => UQVN_N4);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => QI4, A1 => UQVN_N5);
UQVB_B35 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => QI5, A1 => UQVN_N6);
UQVB_B37 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B38 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B39 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => QI6, A1 => UQVN_N7);
UQVB_B40 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => QI7, A1 => UQVN_N8);
UQVB_B41 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N16, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CBD31
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD31 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD31;


ARCHITECTURE lattice_arch OF CBD31 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N3, A1 => UQVN_N7, A2 => UQVN_N8);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => LD);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N7, A1 => CAI, A2 => EN);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => UQVN_N3);
UQVB_B6 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N2, A1 => EN, A2 => CAI);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => LD);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N3);
UQVB_B9 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N1, A1 => UQVN_N6);
UQVB_B10 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N4, A1 => UQVN_N5, A2 => PS);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBD32
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD32 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD32;


ARCHITECTURE lattice_arch OF CBD32 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 QI0, QI1, UQVN_N13, UQVN_N14 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N9, A2 => UQVN_N10);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N9, A1 => CAI, A2 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N13, A1 => CAI, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B8 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N2, A2 => PS);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N9, A2 => UQVN_N10);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => QI0);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => QI1);
UQVB_B12 : AND4
	PORT MAP (Z0 => CAO, A0 => UQVN_N13, A1 => UQVN_N14, A2 => EN, 
	A3 => CAI);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => LD);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B17 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B18 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBD34
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD34;


ARCHITECTURE lattice_arch OF CBD34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, QI0, QI1,
	 QI2, QI3, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N19, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N20, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => D2, A1 => LD);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => D3, A1 => LD);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N23, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN);
UQVB_B12 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N2, A2 => PS);
UQVB_B13 : OR3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => UQVN_N12, A2 => PS);
UQVB_B14 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => UQVN_N16, A2 => PS);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N23, A1 => UQVN_N24, A2 => UQVN_N17, 
	A3 => CAI, A4 => EN);
UQVB_B16 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N23, A1 => UQVN_N24, A2 => UQVN_N25, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI0);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI2);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI3);
UQVB_B22 : AND6
	PORT MAP (Z0 => CAO, A0 => UQVN_N23, A1 => UQVN_N24, A2 => UQVN_N25, 
	A3 => UQVN_N26, A4 => EN, A5 => CAI);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => PS);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B31 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N10, A1 => UQVN_N11);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N14, A1 => UQVN_N15);
END lattice_arch;
-- VHDL netlist for CBD38
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD38;


ARCHITECTURE lattice_arch OF CBD38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 QI0, QI1, QI2, QI3,
	 QI4, QI5, QI6, QI7,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N19, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N20, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => D2, A1 => LD);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => D3, A1 => LD);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N45, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN);
UQVB_B12 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N2, A2 => PS);
UQVB_B13 : OR3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => UQVN_N12, A2 => PS);
UQVB_B14 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => UQVN_N16, A2 => PS);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N17, 
	A3 => CAI, A4 => EN);
UQVB_B16 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => QI0);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => QI1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => QI2);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => QI3);
UQVB_B22 : AND10
	PORT MAP (Z0 => CAO, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N49, A5 => UQVN_N50, A6 => UQVN_N51, 
	A7 => UQVN_N52, A8 => CAI, A9 => EN);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => PS);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B32 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B33 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B35 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B38 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N10, A1 => UQVN_N11);
UQVB_B39 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B40 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => QI4, A1 => UQVN_N25, A2 => UQVN_N37);
UQVB_B41 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => D4, A1 => LD);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => QI5, A1 => UQVN_N25, A2 => UQVN_N37);
UQVB_B43 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => D5, A1 => LD);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => QI6, A1 => UQVN_N25, A2 => UQVN_N37);
UQVB_B45 : AND2
	PORT MAP (Z0 => UQVN_N34, A0 => D6, A1 => LD);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => QI7, A1 => UQVN_N25, A2 => UQVN_N37);
UQVB_B47 : AND2
	PORT MAP (Z0 => UQVN_N40, A0 => D7, A1 => LD);
UQVB_B48 : AND7
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N25, A5 => CAI, A6 => EN);
UQVB_B49 : OR3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N28, A1 => UQVN_N29, A2 => PS);
UQVB_B50 : OR3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N33, A2 => PS);
UQVB_B51 : AND8
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N49, A5 => UQVN_N25, A6 => CAI, 
	A7 => EN);
UQVB_B52 : OR3
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N34, A1 => UQVN_N23, A2 => PS);
UQVB_B53 : AND9
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N49, A5 => UQVN_N50, A6 => UQVN_N25, 
	A7 => CAI, A8 => EN);
UQVB_B54 : AND10
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N45, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N49, A5 => UQVN_N50, A6 => UQVN_N51, 
	A7 => UQVN_N25, A8 => CAI, A9 => EN);
UQVB_B55 : OR3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N24, A2 => PS);
UQVB_B56 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => QI4);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => QI5);
UQVB_B58 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI6);
UQVB_B59 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => QI7);
UQVB_B60 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => PS);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => LD);
UQVB_B62 : LXOR2
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N27, A1 => UQVN_N26);
UQVB_B63 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N41, CLK => CLK, CD => CD);
UQVB_B64 : LXOR2
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N31, A1 => UQVN_N30);
UQVB_B65 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N42, CLK => CLK, CD => CD);
UQVB_B66 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N43, CLK => CLK, CD => CD);
UQVB_B67 : LXOR2
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N35, A1 => UQVN_N36);
UQVB_B68 : LXOR2
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N39, A1 => UQVN_N38);
UQVB_B69 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N44, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CBD41
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD41 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD41;


ARCHITECTURE lattice_arch OF CBD41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N10, CLK => CLK);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => UQVN_N5);
UQVB_B3 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N4, A1 => CAI, A2 => EN);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N7, A2 => UQVN_N9, 
	A3 => UQVN_N8);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => D0, A1 => LD, A2 => UQVN_N9);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N7, A1 => CAI, A2 => EN, 
	A3 => UQVN_N9);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => CS);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => LD);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
UQVB_B10 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N1, A1 => UQVN_N6);
UQVB_B11 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3, A2 => PS);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBD42
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD42 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD42;


ARCHITECTURE lattice_arch OF CBD42 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, QI0, QI1, UQVN_N14,
	 UQVN_N15 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N12, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N13, CLK => CLK);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N4, A2 => PS);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => QI0);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => QI1);
UQVB_B6 : AND4
	PORT MAP (Z0 => CAO, A0 => UQVN_N14, A1 => UQVN_N15, A2 => CAI, 
	A3 => EN);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N9, A2 => UQVN_N11, 
	A3 => UQVN_N10);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => LD, A2 => UQVN_N11);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N9, A1 => CAI, A2 => EN, 
	A3 => UQVN_N11);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N9, A2 => UQVN_N11, 
	A3 => UQVN_N10);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD, A2 => UQVN_N11);
UQVB_B12 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N14, A1 => CAI, A2 => UQVN_N9, 
	A3 => EN, A4 => UQVN_N11);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => CS);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N1, A1 => UQVN_N7);
UQVB_B17 : OR3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => UQVN_N2, A2 => PS);
UQVB_B18 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N3, A1 => UQVN_N8);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => LD);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBD44
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD44;


ARCHITECTURE lattice_arch OF CBD44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, QI0,
	 QI1, QI2, QI3, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N20, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N21, CLK => CLK);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N6, A1 => UQVN_N4, A2 => PS);
UQVB_B4 : OR3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N7, A1 => UQVN_N13, A2 => PS);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N8, A1 => UQVN_N16, A2 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI0);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N19, 
	A3 => UQVN_N18);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => LD, A2 => UQVN_N19);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N17, A1 => CAI, A2 => EN, 
	A3 => UQVN_N19);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N19, 
	A3 => UQVN_N18);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD, A2 => UQVN_N19);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N24, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN, A4 => UQVN_N19);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => D2, A1 => LD, A2 => UQVN_N19);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B18 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N24, A1 => UQVN_N25, A2 => UQVN_N17, 
	A3 => CAI, A4 => EN, A5 => UQVN_N19);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => D3, A1 => LD, A2 => UQVN_N19);
UQVB_B21 : AND7
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N24, A1 => UQVN_N25, A2 => UQVN_N26, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN, A6 => UQVN_N19);
UQVB_B22 : AND6
	PORT MAP (Z0 => CAO, A0 => UQVN_N24, A1 => UQVN_N25, A2 => UQVN_N26, 
	A3 => UQVN_N27, A4 => CAI, A5 => EN);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => CS);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => PS);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B29 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N22, CLK => CLK);
UQVB_B30 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N23, CLK => CLK);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N1, A1 => UQVN_N9);
UQVB_B32 : OR3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N5, A1 => UQVN_N2, A2 => PS);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N3, A1 => UQVN_N10);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N14, A1 => UQVN_N15);
END lattice_arch;
-- VHDL netlist for CBD48
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD48;


ARCHITECTURE lattice_arch OF CBD48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, QI0, QI1,
	 QI2, QI3, QI4, QI5,
	 QI6, QI7, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N20, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N21, CLK => CLK);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N6, A1 => UQVN_N4, A2 => PS);
UQVB_B4 : OR3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N7, A1 => UQVN_N13, A2 => PS);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N8, A1 => UQVN_N16, A2 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => QI0);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => QI1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => QI2);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => QI3);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N19, 
	A3 => UQVN_N18);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => LD, A2 => UQVN_N19);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N17, A1 => CAI, A2 => EN, 
	A3 => UQVN_N19);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N19, 
	A3 => UQVN_N18);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD, A2 => UQVN_N19);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N47, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN, A4 => UQVN_N19);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => D2, A1 => LD, A2 => UQVN_N19);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B18 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N17, 
	A3 => CAI, A4 => EN, A5 => UQVN_N19);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => D3, A1 => LD, A2 => UQVN_N19);
UQVB_B21 : AND7
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN, A6 => UQVN_N19);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => CS);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => PS);
UQVB_B24 : AND10
	PORT MAP (Z0 => CAO, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => UQVN_N50, A4 => UQVN_N51, A5 => UQVN_N52, A6 => UQVN_N53, 
	A7 => UQVN_N54, A8 => CAI, A9 => EN);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B33 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N22, CLK => CLK);
UQVB_B34 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N23, CLK => CLK);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N1, A1 => UQVN_N9);
UQVB_B36 : OR3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N5, A1 => UQVN_N2, A2 => PS);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N3, A1 => UQVN_N10);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B39 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B40 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B41 : OR3
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N30, A1 => UQVN_N31, A2 => PS);
UQVB_B42 : OR3
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N34, A1 => UQVN_N35, A2 => PS);
UQVB_B43 : OR3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N36, A1 => UQVN_N24, A2 => PS);
UQVB_B44 : OR3
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N26, A1 => UQVN_N25, A2 => PS);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI4);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => QI5);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => QI6);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI7);
UQVB_B49 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => QI4, A1 => UQVN_N27, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B50 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => D4, A1 => LD, A2 => UQVN_N40);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => QI5, A1 => UQVN_N27, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => D5, A1 => LD, A2 => UQVN_N40);
UQVB_B53 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => QI6, A1 => UQVN_N27, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B54 : AND3
	PORT MAP (Z0 => UQVN_N36, A0 => D6, A1 => LD, A2 => UQVN_N40);
UQVB_B55 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => UQVN_N27, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B56 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => D7, A1 => LD, A2 => UQVN_N40);
UQVB_B57 : AND11
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => UQVN_N50, A4 => UQVN_N51, A5 => UQVN_N52, A6 => UQVN_N53, 
	A7 => UQVN_N27, A8 => CAI, A9 => EN, A10 => UQVN_N40);
UQVB_B58 : AND10
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => UQVN_N50, A4 => UQVN_N51, A5 => UQVN_N52, A6 => UQVN_N27, 
	A7 => CAI, A8 => EN, A9 => UQVN_N40);
UQVB_B59 : AND9
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => UQVN_N50, A4 => UQVN_N51, A5 => UQVN_N27, A6 => CAI, 
	A7 => EN, A8 => UQVN_N40);
UQVB_B60 : AND8
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => UQVN_N50, A4 => UQVN_N27, A5 => CAI, A6 => EN, 
	A7 => UQVN_N40);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CS);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => PS);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => LD);
UQVB_B64 : LXOR2
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N29, A1 => UQVN_N28);
UQVB_B65 : FD11
	PORT MAP (Q0 => QI4, D0 => UQVN_N43, CLK => CLK);
UQVB_B66 : LXOR2
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N33, A1 => UQVN_N32);
UQVB_B67 : FD11
	PORT MAP (Q0 => QI5, D0 => UQVN_N44, CLK => CLK);
UQVB_B68 : FD11
	PORT MAP (Q0 => QI6, D0 => UQVN_N45, CLK => CLK);
UQVB_B69 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N37, A1 => UQVN_N38);
UQVB_B70 : LXOR2
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N42, A1 => UQVN_N41);
UQVB_B71 : FD11
	PORT MAP (Q0 => QI7, D0 => UQVN_N46, CLK => CLK);
END lattice_arch;
-- VHDL netlist for CBD516
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD516 IS 
    PORT (
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        Q8 : OUT std_logic;
        Q9 : OUT std_logic;
        Q10 : OUT std_logic;
        Q11 : OUT std_logic;
        Q12 : OUT std_logic;
        Q13 : OUT std_logic;
        Q14 : OUT std_logic;
        Q15 : OUT std_logic
    );
END CBD516;


ARCHITECTURE lattice_arch OF CBD516 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, QI0, QI1,
	 QI10, QI11, QI12, QI13,
	 QI14, QI15, QI2, QI3,
	 QI4, QI5, QI6, QI7,
	 QI8, QI9, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


  COMPONENT AND16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND16 use  entity  lat_vhd.AND16(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => EN);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => QI1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => QI2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => QI3);
UQVB_B7 : LXOR2
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => EN);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N5);
UQVB_B9 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI2, A1 => UQVN_N6);
UQVB_B10 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B11 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => UQVN_N7);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q15, A0 => QI15);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q14, A0 => QI14);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q13, A0 => QI13);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q12, A0 => QI12);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q11, A0 => QI11);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q10, A0 => QI10);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q9, A0 => QI9);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q8, A0 => QI8);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B30 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N35, A1 => EN);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N35, A1 => UQVN_N36, A2 => EN);
UQVB_B32 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B33 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B34 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => QI7, A1 => UQVN_N13);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI6, A1 => UQVN_N12);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => QI5, A1 => UQVN_N11);
UQVB_B38 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI4, A1 => UQVN_N14);
UQVB_B39 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => EN);
UQVB_B40 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B41 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => EN);
UQVB_B42 : AND7
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => EN);
UQVB_B43 : AND8
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => EN);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => QI4);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => QI5);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => QI6);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => QI7);
UQVB_B48 : FD21
	PORT MAP (Q0 => QI8, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B49 : FD21
	PORT MAP (Q0 => QI10, D0 => UQVN_N20, CLK => CLK, CD => CD);
UQVB_B50 : FD21
	PORT MAP (Q0 => QI9, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B51 : FD21
	PORT MAP (Q0 => QI11, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B52 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => QI8, A1 => UQVN_N16);
UQVB_B53 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => QI9, A1 => UQVN_N19);
UQVB_B54 : AND9
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => EN);
UQVB_B55 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => QI10, A1 => UQVN_N18);
UQVB_B56 : AND10
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => EN);
UQVB_B57 : AND11
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => UQVN_N49, A10 => EN);
UQVB_B58 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => QI11, A1 => UQVN_N17);
UQVB_B59 : AND12
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => UQVN_N49, A10 => UQVN_N37, 
	A11 => EN);
UQVB_B60 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => QI8);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => QI9);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => QI10);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => QI11);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => QI14);
UQVB_B65 : LXOR2
	PORT MAP (Z0 => UQVN_N26, A0 => QI14, A1 => UQVN_N25);
UQVB_B66 : FD21
	PORT MAP (Q0 => QI15, D0 => UQVN_N32, CLK => CLK, CD => CD);
UQVB_B67 : FD21
	PORT MAP (Q0 => QI13, D0 => UQVN_N28, CLK => CLK, CD => CD);
UQVB_B68 : FD21
	PORT MAP (Q0 => QI12, D0 => UQVN_N29, CLK => CLK, CD => CD);
UQVB_B69 : LXOR2
	PORT MAP (Z0 => UQVN_N28, A0 => QI13, A1 => UQVN_N30);
UQVB_B70 : LXOR2
	PORT MAP (Z0 => UQVN_N29, A0 => QI12, A1 => UQVN_N27);
UQVB_B71 : FD21
	PORT MAP (Q0 => QI14, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => QI15, A1 => UQVN_N24);
UQVB_B73 : AND12
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => UQVN_N49, A10 => UQVN_N37, 
	A11 => UQVN_N38);
UQVB_B74 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N31, A1 => EN);
UQVB_B75 : AND12
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => UQVN_N49, A10 => UQVN_N37, 
	A11 => UQVN_N38);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N33, A1 => UQVN_N39, A2 => EN);
UQVB_B77 : AND12
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => UQVN_N49, A10 => UQVN_N37, 
	A11 => UQVN_N38);
UQVB_B78 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N34, A1 => UQVN_N39, A2 => UQVN_N40, 
	A3 => EN);
UQVB_B79 : AND16
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N35, A1 => UQVN_N36, A2 => UQVN_N42, 
	A3 => UQVN_N43, A4 => UQVN_N44, A5 => UQVN_N45, A6 => UQVN_N46, 
	A7 => UQVN_N47, A8 => UQVN_N48, A9 => UQVN_N49, A10 => UQVN_N37, 
	A11 => UQVN_N38, A12 => UQVN_N39, A13 => UQVN_N40, A14 => UQVN_N41, 
	A15 => EN);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => QI12);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => QI13);
END lattice_arch;
-- VHDL netlist for CBD616
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBD616 IS 
    PORT (
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        Q8 : OUT std_logic;
        Q9 : OUT std_logic;
        Q10 : OUT std_logic;
        Q11 : OUT std_logic;
        Q12 : OUT std_logic;
        Q13 : OUT std_logic;
        Q14 : OUT std_logic;
        Q15 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBD616;


ARCHITECTURE lattice_arch OF CBD616 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, QI0,
	 QI1, QI10, QI11, QI12,
	 QI13, QI14, QI15, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, QI8, QI9, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND16 use  entity  lat_vhd.AND16(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B2 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => EN);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => QI0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => QI1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => QI2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => QI3);
UQVB_B7 : AND2
	PORT MAP (Z0 => CAO, A0 => UQVN_N1, A1 => EN);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => EN);
UQVB_B9 : AND16
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => UQVN_N38, 
	A11 => UQVN_N39, A12 => UQVN_N40, A13 => UQVN_N41, A14 => UQVN_N42, 
	A15 => UQVN_N43);
UQVB_B10 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N6);
UQVB_B11 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI2, A1 => UQVN_N7);
UQVB_B12 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B13 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => UQVN_N8);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q15, A0 => QI15);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q14, A0 => QI14);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q13, A0 => QI13);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q12, A0 => QI12);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q11, A0 => QI11);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q10, A0 => QI10);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q9, A0 => QI9);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q8, A0 => QI8);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B31 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N36, A1 => EN);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N36, A1 => UQVN_N37, A2 => EN);
UQVB_B34 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B35 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B36 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => QI7, A1 => UQVN_N14);
UQVB_B38 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => QI6, A1 => UQVN_N13);
UQVB_B39 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI5, A1 => UQVN_N12);
UQVB_B40 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI4, A1 => UQVN_N15);
UQVB_B41 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => EN);
UQVB_B42 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B43 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => EN);
UQVB_B44 : AND7
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => EN);
UQVB_B45 : AND8
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => EN);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => QI4);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => QI5);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => QI6);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => QI7);
UQVB_B50 : FD21
	PORT MAP (Q0 => QI8, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B51 : FD21
	PORT MAP (Q0 => QI10, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B52 : FD21
	PORT MAP (Q0 => QI9, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B53 : FD21
	PORT MAP (Q0 => QI11, D0 => UQVN_N24, CLK => CLK, CD => CD);
UQVB_B54 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => QI8, A1 => UQVN_N17);
UQVB_B55 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => QI9, A1 => UQVN_N20);
UQVB_B56 : AND9
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => EN);
UQVB_B57 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => QI10, A1 => UQVN_N19);
UQVB_B58 : AND10
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => EN);
UQVB_B59 : AND11
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => EN);
UQVB_B60 : LXOR2
	PORT MAP (Z0 => UQVN_N24, A0 => QI11, A1 => UQVN_N18);
UQVB_B61 : AND12
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => UQVN_N38, 
	A11 => EN);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => QI8);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI9);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => QI10);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => QI11);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => QI14);
UQVB_B67 : LXOR2
	PORT MAP (Z0 => UQVN_N27, A0 => QI14, A1 => UQVN_N26);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => QI15);
UQVB_B69 : FD21
	PORT MAP (Q0 => QI15, D0 => UQVN_N33, CLK => CLK, CD => CD);
UQVB_B70 : FD21
	PORT MAP (Q0 => QI13, D0 => UQVN_N29, CLK => CLK, CD => CD);
UQVB_B71 : FD21
	PORT MAP (Q0 => QI12, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => UQVN_N29, A0 => QI13, A1 => UQVN_N31);
UQVB_B73 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => QI12, A1 => UQVN_N28);
UQVB_B74 : FD21
	PORT MAP (Q0 => QI14, D0 => UQVN_N27, CLK => CLK, CD => CD);
UQVB_B75 : LXOR2
	PORT MAP (Z0 => UQVN_N33, A0 => QI15, A1 => UQVN_N25);
UQVB_B76 : AND12
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => UQVN_N38, 
	A11 => UQVN_N39);
UQVB_B77 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N32, A1 => EN);
UQVB_B78 : AND12
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => UQVN_N38, 
	A11 => UQVN_N39);
UQVB_B79 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N34, A1 => UQVN_N40, A2 => EN);
UQVB_B80 : AND12
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => UQVN_N38, 
	A11 => UQVN_N39);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N35, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => EN);
UQVB_B82 : AND16
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N36, A1 => UQVN_N37, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49, A8 => UQVN_N50, A9 => UQVN_N51, A10 => UQVN_N38, 
	A11 => UQVN_N39, A12 => UQVN_N40, A13 => UQVN_N41, A14 => UQVN_N42, 
	A15 => EN);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => QI12);
UQVB_B84 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => QI13);
END lattice_arch;
-- VHDL netlist for CBU11
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU11 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU11;


ARCHITECTURE lattice_arch OF CBU11 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N1, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B2 : AND2
	PORT MAP (Z0 => CAO, A0 => UQVN_N1, A1 => CAI);
UQVB_B3 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N1);
UQVB_B4 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N1, A1 => CAI);
END lattice_arch;
-- VHDL netlist for CBU12
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU12 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU12;


ARCHITECTURE lattice_arch OF CBU12 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, QI0,
	 QI1 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => CAI);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => CAI);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B7 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for CBU14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU14 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU14;


ARCHITECTURE lattice_arch OF CBU14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, QI0,
	 QI1, QI2, QI3 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B3 : AND5
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => CAI);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => QI1, A2 => CAI);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => CAI);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B11 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B12 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B13 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => CAI);
UQVB_B14 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => QI1, A1 => UQVN_N1);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => UQVN_N6, A0 => QI2, A1 => UQVN_N2);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for CBU18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU18 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU18;


ARCHITECTURE lattice_arch OF CBU18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, QI0,
	 QI1, QI2, QI3, QI4,
	 QI5, QI6, QI7 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => CAI);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => QI1, A2 => CAI);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => CAI);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI);
UQVB_B7 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => CAI);
UQVB_B8 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => CAI);
UQVB_B9 : AND8
	PORT MAP (Z0 => UQVN_N7, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => CAI);
UQVB_B10 : AND9
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => CAI);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B19 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B20 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => QI0, A1 => CAI);
UQVB_B22 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI1, A1 => UQVN_N1);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI2, A1 => UQVN_N2);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => QI3, A1 => UQVN_N3);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => QI4, A1 => UQVN_N4);
UQVB_B26 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B27 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => QI5, A1 => UQVN_N5);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => QI6, A1 => UQVN_N6);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => QI7, A1 => UQVN_N7);
UQVB_B32 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N15, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CBU21
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU21 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU21;


ARCHITECTURE lattice_arch OF CBU21 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B3 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N2, A1 => CAI, A2 => EN);
UQVB_B4 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
UQVB_B5 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N2, A1 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for CBU22
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU22 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU22;


ARCHITECTURE lattice_arch OF CBU22 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 QI0, QI1 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => EN);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI0, A1 => UQVN_N1);
UQVB_B9 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI1, A1 => UQVN_N2);
END lattice_arch;
-- VHDL netlist for CBU24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU24 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU24;


ARCHITECTURE lattice_arch OF CBU24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 QI0, QI1, QI2, QI3 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => EN);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => CAI, A4 => EN);
UQVB_B7 : AND6
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI, A5 => EN);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B12 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B13 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B14 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => UQVN_N1);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => UQVN_N6, A0 => QI1, A1 => UQVN_N2);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => QI2, A1 => UQVN_N3);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => UQVN_N4);
END lattice_arch;
-- VHDL netlist for CBU28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU28 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU28;


ARCHITECTURE lattice_arch OF CBU28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 QI0, QI1, QI2, QI3,
	 QI4, QI5, QI6, QI7 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B3 : AND10
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => CAI, A9 => EN);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => CAI, A1 => EN);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => EN);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => EN);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => CAI, A4 => EN);
UQVB_B8 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI, A5 => EN);
UQVB_B9 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => CAI, A6 => EN);
UQVB_B10 : AND8
	PORT MAP (Z0 => UQVN_N7, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => CAI, 
	A7 => EN);
UQVB_B11 : AND9
	PORT MAP (Z0 => UQVN_N8, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => CAI, A8 => EN);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B20 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B21 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B22 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI0, A1 => UQVN_N1);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI1, A1 => UQVN_N2);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => QI2, A1 => UQVN_N3);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => QI3, A1 => UQVN_N4);
UQVB_B26 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => QI4, A1 => UQVN_N5);
UQVB_B27 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B28 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => QI5, A1 => UQVN_N6);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => QI6, A1 => UQVN_N7);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => QI7, A1 => UQVN_N8);
UQVB_B33 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N16, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CBU31
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU31 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU31;


ARCHITECTURE lattice_arch OF CBU31 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N7, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N7, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => D0, A1 => LD);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => CAI, A2 => EN);
UQVB_B5 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N7, A1 => CAI, A2 => EN);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => LD);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N7);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N1, A1 => UQVN_N4);
UQVB_B9 : OR3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N2, A1 => UQVN_N3, A2 => PS);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBU32
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU32 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU32;


ARCHITECTURE lattice_arch OF CBU32 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 QI0, QI1 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N9, A2 => UQVN_N10);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N9, A1 => CAI, A2 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B8 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N2, A2 => PS);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N9, A2 => UQVN_N10);
UQVB_B10 : AND4
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => EN);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => PS);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B14 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => LD);
END lattice_arch;
-- VHDL netlist for CBU34
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU34;


ARCHITECTURE lattice_arch OF CBU34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, QI0, QI1,
	 QI2, QI3 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N19, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N20, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => D2, A1 => LD);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => D3, A1 => LD);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN);
UQVB_B12 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N2, A2 => PS);
UQVB_B13 : OR3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => UQVN_N12, A2 => PS);
UQVB_B14 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => UQVN_N16, A2 => PS);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => QI0, A1 => QI1, A2 => UQVN_N17, 
	A3 => CAI, A4 => EN);
UQVB_B16 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B18 : AND6
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI, A5 => EN);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => PS);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B24 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B25 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B26 : LXOR2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B27 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B28 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N10, A1 => UQVN_N11);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N14, A1 => UQVN_N15);
END lattice_arch;
-- VHDL netlist for CBU38
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU38;


ARCHITECTURE lattice_arch OF CBU38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 QI0, QI1, QI2, QI3,
	 QI4, QI5, QI6, QI7 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N19, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N20, CLK => CLK, CD => CD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => D2, A1 => LD);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => D3, A1 => LD);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN);
UQVB_B12 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N2, A2 => PS);
UQVB_B13 : OR3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => UQVN_N12, A2 => PS);
UQVB_B14 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => UQVN_N16, A2 => PS);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => QI0, A1 => QI1, A2 => UQVN_N17, 
	A3 => CAI, A4 => EN);
UQVB_B16 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B18 : AND10
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => CAI, A9 => EN);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => PS);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B31 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N10, A1 => UQVN_N11);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B36 : AND10
	PORT MAP (Z0 => UQVN_N25, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => UQVN_N34, A8 => CAI, A9 => EN);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => LD);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => PS);
UQVB_B39 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => QI4, A1 => UQVN_N34, A2 => UQVN_N24);
UQVB_B40 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => QI5, A1 => UQVN_N34, A2 => UQVN_N24);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N44, A0 => QI6, A1 => UQVN_N34, A2 => UQVN_N24);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => UQVN_N34, A2 => UQVN_N24);
UQVB_B43 : AND7
	PORT MAP (Z0 => UQVN_N43, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => UQVN_N34, A5 => CAI, A6 => EN);
UQVB_B44 : AND8
	PORT MAP (Z0 => UQVN_N41, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => UQVN_N34, A6 => CAI, 
	A7 => EN);
UQVB_B45 : AND2
	PORT MAP (Z0 => UQVN_N26, A0 => D5, A1 => LD);
UQVB_B46 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => D4, A1 => LD);
UQVB_B47 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N28, CLK => CLK, CD => CD);
UQVB_B48 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N38, CLK => CLK, CD => CD);
UQVB_B49 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N31, CLK => CLK, CD => CD);
UQVB_B50 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N35, CLK => CLK, CD => CD);
UQVB_B51 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => D6, A1 => LD);
UQVB_B52 : LXOR2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N27, A1 => UQVN_N36);
UQVB_B53 : OR3
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N29, A1 => UQVN_N25, A2 => PS);
UQVB_B54 : AND2
	PORT MAP (Z0 => UQVN_N29, A0 => D7, A1 => LD);
UQVB_B55 : LXOR2
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N44, A1 => UQVN_N37);
UQVB_B56 : OR3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N23, A1 => UQVN_N39, A2 => PS);
UQVB_B57 : LXOR2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N30, A1 => UQVN_N40);
UQVB_B58 : OR3
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N26, A1 => UQVN_N41, A2 => PS);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N33, A1 => UQVN_N42);
UQVB_B60 : OR3
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N32, A1 => UQVN_N43, A2 => PS);
UQVB_B61 : AND9
	PORT MAP (Z0 => UQVN_N39, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => UQVN_N34, 
	A7 => CAI, A8 => EN);
END lattice_arch;
-- VHDL netlist for CBU41
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU41 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU41;


ARCHITECTURE lattice_arch OF CBU41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N9, CLK => CLK);
UQVB_B2 : AND3
	PORT MAP (Z0 => CAO, A0 => UQVN_N2, A1 => CAI, A2 => EN);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => LD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => CS);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD, A2 => UQVN_N7);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N6, A1 => CAI, A2 => EN, 
	A3 => UQVN_N7);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B9 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N7, 
	A3 => UQVN_N8);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBU42
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU42 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU42;


ARCHITECTURE lattice_arch OF CBU42 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, QI0, QI1 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N12, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N13, CLK => CLK);
UQVB_B3 : AND4
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => EN);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => PS);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N9, A1 => CAI, A2 => EN, 
	A3 => UQVN_N10);
UQVB_B10 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N1, A1 => UQVN_N4);
UQVB_B11 : OR3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N2, A1 => UQVN_N3, A2 => PS);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => QI1, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11);
UQVB_B14 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => LD);
UQVB_B17 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => QI0, A1 => CAI, A2 => UQVN_N9, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B18 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N5, A1 => UQVN_N6, A2 => PS);
END lattice_arch;
-- VHDL netlist for CBU44
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU44;


ARCHITECTURE lattice_arch OF CBU44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, QI0,
	 QI1, QI2, QI3 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N20, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N21, CLK => CLK);
UQVB_B3 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => UQVN_N17, A4 => EN, A5 => UQVN_N18);
UQVB_B4 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => UQVN_N16, A2 => PS);
UQVB_B5 : AND7
	PORT MAP (Z0 => UQVN_N16, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN, A6 => UQVN_N18);
UQVB_B6 : AND6
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI, A5 => EN);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => CS);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => PS);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B13 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N22, CLK => CLK);
UQVB_B14 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N23, CLK => CLK);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD, A2 => UQVN_N18);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => EN, 
	A3 => UQVN_N18);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B18 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B20 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD, A2 => UQVN_N18);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D2, A1 => LD, A2 => UQVN_N18);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B26 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B27 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => D3, A1 => LD, A2 => UQVN_N18);
UQVB_B29 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B30 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI0, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN, A4 => UQVN_N18);
UQVB_B31 : OR3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N6, A1 => UQVN_N7, A2 => PS);
UQVB_B32 : OR3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N10, A1 => UQVN_N2, A2 => PS);
END lattice_arch;
-- VHDL netlist for CBU48
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU48;


ARCHITECTURE lattice_arch OF CBU48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, QI0, QI1,
	 QI2, QI3, QI4, QI5,
	 QI6, QI7 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N20, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N21, CLK => CLK);
UQVB_B3 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => UQVN_N17, A4 => EN, A5 => UQVN_N18);
UQVB_B4 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => UQVN_N16, A2 => PS);
UQVB_B5 : AND7
	PORT MAP (Z0 => UQVN_N16, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N17, A4 => CAI, A5 => EN, A6 => UQVN_N18);
UQVB_B6 : AND10
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => CAI, A9 => EN);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => CS);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => PS);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B17 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N22, CLK => CLK);
UQVB_B18 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N23, CLK => CLK);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => LD, A2 => UQVN_N18);
UQVB_B20 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => EN, 
	A3 => UQVN_N18);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N1, A1 => UQVN_N5);
UQVB_B22 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N3, A1 => UQVN_N4, A2 => PS);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B24 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => QI1, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => D1, A1 => LD, A2 => UQVN_N18);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D2, A1 => LD, A2 => UQVN_N18);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B30 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => QI2, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => D3, A1 => LD, A2 => UQVN_N18);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => UQVN_N17, A2 => UQVN_N18, 
	A3 => UQVN_N19);
UQVB_B34 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI0, A1 => CAI, A2 => UQVN_N17, 
	A3 => EN, A4 => UQVN_N18);
UQVB_B35 : OR3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N6, A1 => UQVN_N7, A2 => PS);
UQVB_B36 : OR3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N10, A1 => UQVN_N2, A2 => PS);
UQVB_B37 : AND8
	PORT MAP (Z0 => UQVN_N29, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => UQVN_N25, A5 => CAI, A6 => EN, 
	A7 => UQVN_N38);
UQVB_B38 : AND9
	PORT MAP (Z0 => UQVN_N33, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => UQVN_N25, A6 => CAI, 
	A7 => EN, A8 => UQVN_N38);
UQVB_B39 : AND10
	PORT MAP (Z0 => UQVN_N34, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => UQVN_N25, 
	A7 => CAI, A8 => EN, A9 => UQVN_N38);
UQVB_B40 : AND11
	PORT MAP (Z0 => UQVN_N24, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => UQVN_N25, A8 => CAI, A9 => EN, A10 => UQVN_N38);
UQVB_B41 : OR3
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N42, A1 => UQVN_N24, A2 => PS);
UQVB_B42 : OR3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N28, A1 => UQVN_N29, A2 => PS);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => CS);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => LD);
UQVB_B45 : LXOR2
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N27, A1 => UQVN_N26);
UQVB_B46 : FD11
	PORT MAP (Q0 => QI4, D0 => UQVN_N43, CLK => CLK);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => D4, A1 => LD, A2 => UQVN_N38);
UQVB_B48 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => QI4, A1 => UQVN_N25, A2 => UQVN_N38, 
	A3 => UQVN_N39);
UQVB_B49 : LXOR2
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N31, A1 => UQVN_N30);
UQVB_B50 : FD11
	PORT MAP (Q0 => QI5, D0 => UQVN_N44, CLK => CLK);
UQVB_B51 : OR3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N33, A2 => PS);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N32, A0 => D5, A1 => LD, A2 => UQVN_N38);
UQVB_B53 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => QI5, A1 => UQVN_N25, A2 => UQVN_N38, 
	A3 => UQVN_N39);
UQVB_B54 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => D6, A1 => LD, A2 => UQVN_N38);
UQVB_B55 : OR3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N35, A1 => UQVN_N34, A2 => PS);
UQVB_B56 : FD11
	PORT MAP (Q0 => QI6, D0 => UQVN_N45, CLK => CLK);
UQVB_B57 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N36, A1 => UQVN_N37);
UQVB_B58 : AND4
	PORT MAP (Z0 => UQVN_N36, A0 => QI6, A1 => UQVN_N25, A2 => UQVN_N38, 
	A3 => UQVN_N39);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N41, A1 => UQVN_N40);
UQVB_B60 : FD11
	PORT MAP (Q0 => QI7, D0 => UQVN_N46, CLK => CLK);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N42, A0 => D7, A1 => LD, A2 => UQVN_N38);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => UQVN_N25, A2 => UQVN_N38, 
	A3 => UQVN_N39);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => PS);
END lattice_arch;
-- VHDL netlist for CBU516
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU516 IS 
    PORT (
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        Q8 : OUT std_logic;
        Q9 : OUT std_logic;
        Q10 : OUT std_logic;
        Q11 : OUT std_logic;
        Q12 : OUT std_logic;
        Q13 : OUT std_logic;
        Q14 : OUT std_logic;
        Q15 : OUT std_logic
    );
END CBU516;


ARCHITECTURE lattice_arch OF CBU516 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, QI0, QI1,
	 QI10, QI11, QI12, QI13,
	 QI14, QI15, QI2, QI3,
	 QI4, QI5, QI6, QI7,
	 QI8, QI9 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


  COMPONENT AND16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND16 use  entity  lat_vhd.AND16(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => EN);
UQVB_B3 : LXOR2
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => EN);
UQVB_B4 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N5);
UQVB_B5 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI2, A1 => UQVN_N6);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q15, A0 => QI15);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q14, A0 => QI14);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q13, A0 => QI13);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q12, A0 => QI12);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q11, A0 => QI11);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q10, A0 => QI10);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q9, A0 => QI9);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q8, A0 => QI8);
UQVB_B14 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => UQVN_N7);
UQVB_B24 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B25 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => EN);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => QI0, A1 => QI1, A2 => EN);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => QI7, A1 => UQVN_N13);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI6, A1 => UQVN_N12);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => QI5, A1 => UQVN_N11);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI4, A1 => UQVN_N14);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => EN);
UQVB_B36 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B37 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => EN);
UQVB_B38 : AND7
	PORT MAP (Z0 => UQVN_N12, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => EN);
UQVB_B39 : AND8
	PORT MAP (Z0 => UQVN_N13, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => EN);
UQVB_B40 : FD21
	PORT MAP (Q0 => QI8, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B41 : FD21
	PORT MAP (Q0 => QI10, D0 => UQVN_N20, CLK => CLK, CD => CD);
UQVB_B42 : FD21
	PORT MAP (Q0 => QI9, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B43 : FD21
	PORT MAP (Q0 => QI11, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B44 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => QI8, A1 => UQVN_N16);
UQVB_B45 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => QI9, A1 => UQVN_N19);
UQVB_B46 : AND9
	PORT MAP (Z0 => UQVN_N16, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => EN);
UQVB_B47 : LXOR2
	PORT MAP (Z0 => UQVN_N20, A0 => QI10, A1 => UQVN_N18);
UQVB_B48 : AND10
	PORT MAP (Z0 => UQVN_N19, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => EN);
UQVB_B49 : AND11
	PORT MAP (Z0 => UQVN_N18, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => EN);
UQVB_B50 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => QI11, A1 => UQVN_N17);
UQVB_B51 : AND12
	PORT MAP (Z0 => UQVN_N17, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => EN);
UQVB_B52 : LXOR2
	PORT MAP (Z0 => UQVN_N26, A0 => QI14, A1 => UQVN_N25);
UQVB_B53 : FD21
	PORT MAP (Q0 => QI15, D0 => UQVN_N32, CLK => CLK, CD => CD);
UQVB_B54 : FD21
	PORT MAP (Q0 => QI13, D0 => UQVN_N28, CLK => CLK, CD => CD);
UQVB_B55 : FD21
	PORT MAP (Q0 => QI12, D0 => UQVN_N29, CLK => CLK, CD => CD);
UQVB_B56 : LXOR2
	PORT MAP (Z0 => UQVN_N28, A0 => QI13, A1 => UQVN_N30);
UQVB_B57 : LXOR2
	PORT MAP (Z0 => UQVN_N29, A0 => QI12, A1 => UQVN_N27);
UQVB_B58 : FD21
	PORT MAP (Q0 => QI14, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => QI15, A1 => UQVN_N24);
UQVB_B60 : AND12
	PORT MAP (Z0 => UQVN_N31, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11);
UQVB_B61 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N31, A1 => EN);
UQVB_B62 : AND12
	PORT MAP (Z0 => UQVN_N33, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11);
UQVB_B63 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N33, A1 => QI12, A2 => EN);
UQVB_B64 : AND12
	PORT MAP (Z0 => UQVN_N34, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11);
UQVB_B65 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N34, A1 => QI12, A2 => QI13, 
	A3 => EN);
UQVB_B66 : AND16
	PORT MAP (Z0 => UQVN_N24, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => QI13, A14 => QI14, 
	A15 => EN);
END lattice_arch;
-- VHDL netlist for CBU616
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU616 IS 
    PORT (
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        Q8 : OUT std_logic;
        Q9 : OUT std_logic;
        Q10 : OUT std_logic;
        Q11 : OUT std_logic;
        Q12 : OUT std_logic;
        Q13 : OUT std_logic;
        Q14 : OUT std_logic;
        Q15 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBU616;


ARCHITECTURE lattice_arch OF CBU616 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, QI0,
	 QI1, QI10, QI11, QI12,
	 QI13, QI14, QI15, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, QI8, QI9 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND16 use  entity  lat_vhd.AND16(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B2 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => EN);
UQVB_B3 : AND16
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => QI13, A14 => QI14, 
	A15 => QI15);
UQVB_B4 : AND2
	PORT MAP (Z0 => CAO, A0 => UQVN_N1, A1 => EN);
UQVB_B5 : LXOR2
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => EN);
UQVB_B6 : LXOR2
	PORT MAP (Z0 => UQVN_N3, A0 => QI1, A1 => UQVN_N6);
UQVB_B7 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => QI2, A1 => UQVN_N7);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q15, A0 => QI15);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q14, A0 => QI14);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q13, A0 => QI13);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q12, A0 => QI12);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q11, A0 => QI11);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q10, A0 => QI10);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q9, A0 => QI9);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q8, A0 => QI8);
UQVB_B16 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => UQVN_N8);
UQVB_B26 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B27 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => QI0, A1 => EN);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => QI0, A1 => QI1, A2 => EN);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B31 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B32 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => QI7, A1 => UQVN_N14);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => QI6, A1 => UQVN_N13);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => QI5, A1 => UQVN_N12);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => QI4, A1 => UQVN_N15);
UQVB_B37 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => EN);
UQVB_B38 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B39 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => EN);
UQVB_B40 : AND7
	PORT MAP (Z0 => UQVN_N13, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => EN);
UQVB_B41 : AND8
	PORT MAP (Z0 => UQVN_N14, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => EN);
UQVB_B42 : FD21
	PORT MAP (Q0 => QI8, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B43 : FD21
	PORT MAP (Q0 => QI10, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B44 : FD21
	PORT MAP (Q0 => QI9, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B45 : FD21
	PORT MAP (Q0 => QI11, D0 => UQVN_N24, CLK => CLK, CD => CD);
UQVB_B46 : LXOR2
	PORT MAP (Z0 => UQVN_N22, A0 => QI8, A1 => UQVN_N17);
UQVB_B47 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => QI9, A1 => UQVN_N20);
UQVB_B48 : AND9
	PORT MAP (Z0 => UQVN_N17, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => EN);
UQVB_B49 : LXOR2
	PORT MAP (Z0 => UQVN_N21, A0 => QI10, A1 => UQVN_N19);
UQVB_B50 : AND10
	PORT MAP (Z0 => UQVN_N20, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => EN);
UQVB_B51 : AND11
	PORT MAP (Z0 => UQVN_N19, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => EN);
UQVB_B52 : LXOR2
	PORT MAP (Z0 => UQVN_N24, A0 => QI11, A1 => UQVN_N18);
UQVB_B53 : AND12
	PORT MAP (Z0 => UQVN_N18, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => EN);
UQVB_B54 : LXOR2
	PORT MAP (Z0 => UQVN_N27, A0 => QI14, A1 => UQVN_N26);
UQVB_B55 : FD21
	PORT MAP (Q0 => QI15, D0 => UQVN_N33, CLK => CLK, CD => CD);
UQVB_B56 : FD21
	PORT MAP (Q0 => QI13, D0 => UQVN_N29, CLK => CLK, CD => CD);
UQVB_B57 : FD21
	PORT MAP (Q0 => QI12, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B58 : LXOR2
	PORT MAP (Z0 => UQVN_N29, A0 => QI13, A1 => UQVN_N31);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => QI12, A1 => UQVN_N28);
UQVB_B60 : FD21
	PORT MAP (Q0 => QI14, D0 => UQVN_N27, CLK => CLK, CD => CD);
UQVB_B61 : LXOR2
	PORT MAP (Z0 => UQVN_N33, A0 => QI15, A1 => UQVN_N25);
UQVB_B62 : AND12
	PORT MAP (Z0 => UQVN_N32, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11);
UQVB_B63 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N32, A1 => EN);
UQVB_B64 : AND12
	PORT MAP (Z0 => UQVN_N34, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11);
UQVB_B65 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N34, A1 => QI12, A2 => EN);
UQVB_B66 : AND12
	PORT MAP (Z0 => UQVN_N35, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11);
UQVB_B67 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N35, A1 => QI12, A2 => QI13, 
	A3 => EN);
UQVB_B68 : AND16
	PORT MAP (Z0 => UQVN_N25, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => QI13, A14 => QI14, 
	A15 => EN);
END lattice_arch;
-- VHDL netlist for CBU716
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBU716 IS 
    PORT (
        CAI : IN std_logic;
        CD : IN std_logic;
        CLK : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        D10 : IN std_logic;
        D11 : IN std_logic;
        D12 : IN std_logic;
        D13 : IN std_logic;
        D14 : IN std_logic;
        D15 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        D8 : IN std_logic;
        D9 : IN std_logic;
        EN : IN std_logic;
        LD : IN std_logic;
        CAO : OUT std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q10 : OUT std_logic;
        Q11 : OUT std_logic;
        Q12 : OUT std_logic;
        Q13 : OUT std_logic;
        Q14 : OUT std_logic;
        Q15 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        Q8 : OUT std_logic;
        Q9 : OUT std_logic
    );
END CBU716;


ARCHITECTURE lattice_arch OF CBU716 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, QI0, QI1, QI10,
	 QI11, QI12, QI13, QI14,
	 QI15, QI2, QI3, QI4,
	 QI5, QI6, QI7, QI8,
	 QI9 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND18
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        A16 : IN std_logic;
        A17 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND18 use  entity  lat_vhd.AND18(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


  COMPONENT AND13
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND13 use  entity  lat_vhd.AND13(lattice_arch);


  COMPONENT AND14
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND14 use  entity  lat_vhd.AND14(lattice_arch);


  COMPONENT AND15
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND15 use  entity  lat_vhd.AND15(lattice_arch);


  COMPONENT AND16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND16 use  entity  lat_vhd.AND16(lattice_arch);


  COMPONENT AND17
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        A16 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND17 use  entity  lat_vhd.AND17(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N24, CLK => CLK, CD => CD);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => D0, A1 => LD);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N22, A1 => CAI, A2 => EN);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => D1, A1 => LD);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => D2, A1 => LD);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => D3, A1 => LD);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => CAI, A2 => UQVN_N22, 
	A3 => EN);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N17, A0 => QI0, A1 => QI1, A2 => UQVN_N22, 
	A3 => CAI, A4 => EN);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N21, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N22, A4 => CAI, A5 => EN);
UQVB_B11 : AND18
	PORT MAP (Z0 => CAO, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => QI13, A14 => QI14, 
	A15 => QI15, A16 => CAI, A17 => EN);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N22);
UQVB_B13 : OR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q15, A0 => QI15);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q11, A0 => QI11);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q9, A0 => QI9);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q8, A0 => QI8);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q14, A0 => QI14);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q13, A0 => QI13);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q12, A0 => QI12);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q10, A0 => QI10);
UQVB_B30 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => QI1, A1 => UQVN_N22);
UQVB_B31 : OR2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N11, A1 => UQVN_N2);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => QI2, A1 => UQVN_N22);
UQVB_B33 : OR2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N14, A1 => UQVN_N17);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => QI3, A1 => UQVN_N22);
UQVB_B35 : OR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N18, A1 => UQVN_N21);
UQVB_B36 : OR2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N3, A1 => UQVN_N5);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => QI4, A1 => UQVN_N22);
UQVB_B38 : LXOR2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N6, A1 => UQVN_N7);
UQVB_B39 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D4, A1 => LD);
UQVB_B41 : AND7
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => UQVN_N22, A5 => CAI, A6 => EN);
UQVB_B42 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N25, CLK => CLK, CD => CD);
UQVB_B43 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B44 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N1, A1 => UQVN_N10);
UQVB_B45 : LXOR2
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N12, A1 => UQVN_N13);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => LD);
UQVB_B47 : LXOR2
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N15, A1 => UQVN_N16);
UQVB_B48 : LXOR2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N19, A1 => UQVN_N20);
UQVB_B49 : AND10
	PORT MAP (Z0 => UQVN_N33, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => UQVN_N40, A8 => CAI, A9 => EN);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => LD);
UQVB_B51 : AND2
	PORT MAP (Z0 => UQVN_N38, A0 => QI5, A1 => UQVN_N40);
UQVB_B52 : OR2
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N34, A1 => UQVN_N46);
UQVB_B53 : AND2
	PORT MAP (Z0 => UQVN_N47, A0 => QI6, A1 => UQVN_N40);
UQVB_B54 : OR2
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N27, A1 => UQVN_N44);
UQVB_B55 : AND2
	PORT MAP (Z0 => UQVN_N35, A0 => QI7, A1 => UQVN_N40);
UQVB_B56 : OR2
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N37, A1 => UQVN_N33);
UQVB_B57 : OR2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N28, A1 => UQVN_N32);
UQVB_B58 : AND2
	PORT MAP (Z0 => UQVN_N30, A0 => QI8, A1 => UQVN_N40);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N30, A1 => UQVN_N31);
UQVB_B60 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => D8, A1 => LD);
UQVB_B61 : FD21
	PORT MAP (Q0 => QI8, D0 => UQVN_N29, CLK => CLK, CD => CD);
UQVB_B62 : AND11
	PORT MAP (Z0 => UQVN_N32, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => UQVN_N40, A9 => CAI, A10 => EN);
UQVB_B63 : AND8
	PORT MAP (Z0 => UQVN_N46, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => UQVN_N40, A6 => CAI, 
	A7 => EN);
UQVB_B64 : AND2
	PORT MAP (Z0 => UQVN_N34, A0 => D5, A1 => LD);
UQVB_B65 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N36, CLK => CLK, CD => CD);
UQVB_B66 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N43, CLK => CLK, CD => CD);
UQVB_B67 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N39, CLK => CLK, CD => CD);
UQVB_B68 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => D6, A1 => LD);
UQVB_B69 : LXOR2
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N35, A1 => UQVN_N41);
UQVB_B70 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => D7, A1 => LD);
UQVB_B71 : LXOR2
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N47, A1 => UQVN_N42);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N38, A1 => UQVN_N45);
UQVB_B73 : AND9
	PORT MAP (Z0 => UQVN_N44, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => UQVN_N40, 
	A7 => CAI, A8 => EN);
UQVB_B74 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => LD);
UQVB_B75 : AND2
	PORT MAP (Z0 => UQVN_N54, A0 => QI9, A1 => UQVN_N56);
UQVB_B76 : OR2
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N50, A1 => UQVN_N62);
UQVB_B77 : AND2
	PORT MAP (Z0 => UQVN_N63, A0 => QI10, A1 => UQVN_N56);
UQVB_B78 : OR2
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N48, A1 => UQVN_N60);
UQVB_B79 : AND2
	PORT MAP (Z0 => UQVN_N51, A0 => QI11, A1 => UQVN_N56);
UQVB_B80 : OR2
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N53, A1 => UQVN_N49);
UQVB_B81 : AND12
	PORT MAP (Z0 => UQVN_N62, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => UQVN_N56, A10 => CAI, 
	A11 => EN);
UQVB_B82 : AND13
	PORT MAP (Z0 => UQVN_N60, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => UQVN_N56, 
	A11 => CAI, A12 => EN);
UQVB_B83 : AND14
	PORT MAP (Z0 => UQVN_N49, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => UQVN_N56, A12 => CAI, A13 => EN);
UQVB_B84 : AND2
	PORT MAP (Z0 => UQVN_N50, A0 => D9, A1 => LD);
UQVB_B85 : FD21
	PORT MAP (Q0 => QI11, D0 => UQVN_N52, CLK => CLK, CD => CD);
UQVB_B86 : FD21
	PORT MAP (Q0 => QI10, D0 => UQVN_N59, CLK => CLK, CD => CD);
UQVB_B87 : FD21
	PORT MAP (Q0 => QI9, D0 => UQVN_N55, CLK => CLK, CD => CD);
UQVB_B88 : AND2
	PORT MAP (Z0 => UQVN_N48, A0 => D10, A1 => LD);
UQVB_B89 : LXOR2
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N51, A1 => UQVN_N57);
UQVB_B90 : AND2
	PORT MAP (Z0 => UQVN_N53, A0 => D11, A1 => LD);
UQVB_B91 : LXOR2
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N63, A1 => UQVN_N58);
UQVB_B92 : LXOR2
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N54, A1 => UQVN_N61);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N64, A0 => LD);
UQVB_B94 : AND2
	PORT MAP (Z0 => UQVN_N69, A0 => QI12, A1 => UQVN_N64);
UQVB_B95 : OR2
	PORT MAP (Z0 => UQVN_N73, A0 => UQVN_N68, A1 => UQVN_N74);
UQVB_B96 : AND2
	PORT MAP (Z0 => UQVN_N66, A0 => QI13, A1 => UQVN_N64);
UQVB_B97 : OR2
	PORT MAP (Z0 => UQVN_N71, A0 => UQVN_N65, A1 => UQVN_N72);
UQVB_B98 : AND15
	PORT MAP (Z0 => UQVN_N74, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => UQVN_N64, A13 => CAI, A14 => EN);
UQVB_B99 : AND16
	PORT MAP (Z0 => UQVN_N72, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => UQVN_N64, A14 => CAI, 
	A15 => EN);
UQVB_B100 : AND2
	PORT MAP (Z0 => UQVN_N65, A0 => D13, A1 => LD);
UQVB_B101 : AND2
	PORT MAP (Z0 => UQVN_N68, A0 => D12, A1 => LD);
UQVB_B102 : FD21
	PORT MAP (Q0 => QI13, D0 => UQVN_N67, CLK => CLK, CD => CD);
UQVB_B103 : FD21
	PORT MAP (Q0 => QI12, D0 => UQVN_N70, CLK => CLK, CD => CD);
UQVB_B104 : LXOR2
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N66, A1 => UQVN_N71);
UQVB_B105 : LXOR2
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N69, A1 => UQVN_N73);
UQVB_B106 : INV
	PORT MAP (ZN0 => UQVN_N80, A0 => LD);
UQVB_B107 : AND2
	PORT MAP (Z0 => UQVN_N85, A0 => QI14, A1 => UQVN_N80);
UQVB_B108 : OR2
	PORT MAP (Z0 => UQVN_N82, A0 => UQVN_N75, A1 => UQVN_N84);
UQVB_B109 : AND2
	PORT MAP (Z0 => UQVN_N77, A0 => QI15, A1 => UQVN_N80);
UQVB_B110 : OR2
	PORT MAP (Z0 => UQVN_N81, A0 => UQVN_N79, A1 => UQVN_N76);
UQVB_B111 : AND17
	PORT MAP (Z0 => UQVN_N84, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => QI13, A14 => UQVN_N80, 
	A15 => CAI, A16 => EN);
UQVB_B112 : AND18
	PORT MAP (Z0 => UQVN_N76, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => QI8, A9 => QI9, A10 => QI10, 
	A11 => QI11, A12 => QI12, A13 => QI13, A14 => QI14, 
	A15 => UQVN_N80, A16 => CAI, A17 => EN);
UQVB_B113 : FD21
	PORT MAP (Q0 => QI15, D0 => UQVN_N78, CLK => CLK, CD => CD);
UQVB_B114 : FD21
	PORT MAP (Q0 => QI14, D0 => UQVN_N83, CLK => CLK, CD => CD);
UQVB_B115 : AND2
	PORT MAP (Z0 => UQVN_N75, A0 => D14, A1 => LD);
UQVB_B116 : LXOR2
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N77, A1 => UQVN_N81);
UQVB_B117 : AND2
	PORT MAP (Z0 => UQVN_N79, A0 => D15, A1 => LD);
UQVB_B118 : LXOR2
	PORT MAP (Z0 => UQVN_N83, A0 => UQVN_N85, A1 => UQVN_N82);
END lattice_arch;
-- VHDL netlist for CBUD1
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBUD1 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBUD1;


ARCHITECTURE lattice_arch OF CBUD1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UP : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N8, A1 => UQVN_N10, A2 => PS);
UQVB_B2 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N1, A1 => UQVN_N9);
UQVB_B3 : OR2
	PORT MAP (Z0 => CAO, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N3, A1 => CAI, A2 => EN, 
	A3 => DNUP);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N2, A1 => CAI, A2 => EN, 
	A3 => UP);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => UQVN_N2);
UQVB_B7 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => PS);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => UQVN_N5, A2 => UQVN_N4, 
	A3 => UQVN_N6);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => D0, A1 => LD, A2 => UQVN_N4);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N5, A1 => CAI, A2 => EN, 
	A3 => UQVN_N4);
UQVB_B12 : INV
	PORT MAP (ZN0 => UP, A0 => DNUP);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => LD);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
END lattice_arch;
-- VHDL netlist for CBUD2
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBUD2 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBUD2;


ARCHITECTURE lattice_arch OF CBUD2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 QI0, QI1, UP, UQVN_N17,
	 UQVN_N18 : std_logic;


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N1, A1 => UQVN_N9);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N12, A1 => UQVN_N14, A2 => PS);
UQVB_B3 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N2, A1 => UQVN_N13);
UQVB_B4 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N3, A1 => UQVN_N5, A2 => UQVN_N4, 
	A3 => PS);
UQVB_B5 : OR2
	PORT MAP (Z0 => CAO, A0 => UQVN_N15, A1 => UQVN_N16);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N17, A1 => UQVN_N18, A2 => CAI, 
	A3 => EN, A4 => DNUP);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => QI0);
UQVB_B8 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B9 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => QI1);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI0, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N8);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI1, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N8);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => D0, A1 => LD, A2 => UQVN_N6);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N7, A1 => CAI, A2 => EN, 
	A3 => UQVN_N6);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD, A2 => UQVN_N6);
UQVB_B16 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI0, A1 => CAI, A2 => UQVN_N7, 
	A3 => EN, A4 => UQVN_N6, A5 => UP);
UQVB_B17 : AND6
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => CAI, A2 => UQVN_N7, 
	A3 => EN, A4 => UQVN_N6, A5 => DNUP);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => LD);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => CS);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => PS);
UQVB_B21 : INV
	PORT MAP (ZN0 => UP, A0 => DNUP);
UQVB_B22 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => QI0, A1 => QI1, A2 => CAI, 
	A3 => EN, A4 => UP);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
END lattice_arch;
-- VHDL netlist for CBUD4
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBUD4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBUD4;


ARCHITECTURE lattice_arch OF CBUD4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, QI0,
	 QI1, QI2, QI3, UP,
	 UQVN_N32, UQVN_N33, UQVN_N34, UQVN_N35 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B3 : OR2
	PORT MAP (Z0 => CAO, A0 => UQVN_N4, A1 => UQVN_N3);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CS);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UP, A0 => DNUP);
UQVB_B7 : AND7
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N32, A1 => UQVN_N33, A2 => UQVN_N34, 
	A3 => UQVN_N35, A4 => CAI, A5 => EN, A6 => DNUP);
UQVB_B8 : AND7
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => CAI, A5 => EN, A6 => UP);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => LD, A2 => UQVN_N2);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N12, A1 => CAI, A2 => EN, 
	A3 => UQVN_N2);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N1, A1 => UQVN_N7);
UQVB_B16 : OR3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => UQVN_N6, A2 => PS);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N12, A2 => UQVN_N2, 
	A3 => UQVN_N14);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => QI1, A1 => UQVN_N12, A2 => UQVN_N2, 
	A3 => UQVN_N14);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N10, A1 => UQVN_N11);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => D1, A1 => LD, A2 => UQVN_N2);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => LD);
UQVB_B22 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => QI0, A1 => CAI, A2 => UQVN_N12, 
	A3 => EN, A4 => UQVN_N2, A5 => UP);
UQVB_B23 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N32, A1 => CAI, A2 => UQVN_N12, 
	A3 => EN, A4 => UQVN_N2, A5 => DNUP);
UQVB_B24 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N13, 
	A3 => PS);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => QI0);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => QI1);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => CS);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => PS);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N31, CLK => CLK, CD => CD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => LD);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => D2, A1 => LD, A2 => UQVN_N17);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N19, A1 => UQVN_N20);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N26, A2 => UQVN_N17, 
	A3 => UQVN_N29);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N23, A1 => UQVN_N24);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D3, A1 => LD, A2 => UQVN_N17);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => UQVN_N26, A2 => UQVN_N17, 
	A3 => UQVN_N29);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => QI2);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => QI3);
UQVB_B40 : AND7
	PORT MAP (Z0 => UQVN_N21, A0 => QI0, A1 => QI1, A2 => UQVN_N26, 
	A3 => CAI, A4 => EN, A5 => UQVN_N17, A6 => UP);
UQVB_B41 : AND7
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N32, A1 => UQVN_N33, A2 => UQVN_N26, 
	A3 => CAI, A4 => EN, A5 => UQVN_N17, A6 => DNUP);
UQVB_B42 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N18, A1 => UQVN_N21, A2 => UQVN_N27, 
	A3 => PS);
UQVB_B43 : AND8
	PORT MAP (Z0 => UQVN_N25, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N26, A4 => CAI, A5 => EN, A6 => UQVN_N17, 
	A7 => UP);
UQVB_B44 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N32, A1 => UQVN_N33, A2 => UQVN_N34, 
	A3 => UQVN_N26, A4 => CAI, A5 => EN, A6 => UQVN_N17, 
	A7 => DNUP);
UQVB_B45 : OR4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N22, A1 => UQVN_N25, A2 => UQVN_N28, 
	A3 => PS);
END lattice_arch;
-- VHDL netlist for CBUD8
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CBUD8 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CBUD8;


ARCHITECTURE lattice_arch OF CBUD8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, QI0, QI1, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, UP, UQVN_N62, UQVN_N63,
	 UQVN_N64, UQVN_N65, UQVN_N66, UQVN_N67,
	 UQVN_N68, UQVN_N69 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B3 : OR2
	PORT MAP (Z0 => CAO, A0 => UQVN_N4, A1 => UQVN_N3);
UQVB_B4 : AND11
	PORT MAP (Z0 => UQVN_N4, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => QI7, A8 => CAI, A9 => EN, A10 => UP);
UQVB_B5 : AND11
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N65, A4 => UQVN_N66, A5 => UQVN_N67, A6 => UQVN_N68, 
	A7 => UQVN_N69, A8 => CAI, A9 => EN, A10 => DNUP);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CS);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => PS);
UQVB_B8 : INV
	PORT MAP (ZN0 => UP, A0 => DNUP);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => LD, A2 => UQVN_N2);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N12, A1 => CAI, A2 => EN, 
	A3 => UQVN_N2);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N1, A1 => UQVN_N7);
UQVB_B20 : OR3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => UQVN_N6, A2 => PS);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => QI0, A1 => UQVN_N12, A2 => UQVN_N2, 
	A3 => UQVN_N14);
UQVB_B22 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => QI1, A1 => UQVN_N12, A2 => UQVN_N2, 
	A3 => UQVN_N14);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N10, A1 => UQVN_N11);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => D1, A1 => LD, A2 => UQVN_N2);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => LD);
UQVB_B26 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => QI0, A1 => CAI, A2 => UQVN_N12, 
	A3 => EN, A4 => UQVN_N2, A5 => UP);
UQVB_B27 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N62, A1 => CAI, A2 => UQVN_N12, 
	A3 => EN, A4 => UQVN_N2, A5 => DNUP);
UQVB_B28 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N13, 
	A3 => PS);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => QI0);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N63, A0 => QI1);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => CS);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => PS);
UQVB_B33 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B34 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N31, CLK => CLK, CD => CD);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => LD);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => D2, A1 => LD, A2 => UQVN_N17);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N19, A1 => UQVN_N20);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N26, A2 => UQVN_N17, 
	A3 => UQVN_N29);
UQVB_B39 : LXOR2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N23, A1 => UQVN_N24);
UQVB_B40 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D3, A1 => LD, A2 => UQVN_N17);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => UQVN_N26, A2 => UQVN_N17, 
	A3 => UQVN_N29);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N64, A0 => QI2);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => QI3);
UQVB_B44 : AND7
	PORT MAP (Z0 => UQVN_N21, A0 => QI0, A1 => QI1, A2 => UQVN_N26, 
	A3 => CAI, A4 => EN, A5 => UQVN_N17, A6 => UP);
UQVB_B45 : AND7
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N26, 
	A3 => CAI, A4 => EN, A5 => UQVN_N17, A6 => DNUP);
UQVB_B46 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N18, A1 => UQVN_N21, A2 => UQVN_N27, 
	A3 => PS);
UQVB_B47 : AND8
	PORT MAP (Z0 => UQVN_N25, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => UQVN_N26, A4 => CAI, A5 => EN, A6 => UQVN_N17, 
	A7 => UP);
UQVB_B48 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N26, A4 => CAI, A5 => EN, A6 => UQVN_N17, 
	A7 => DNUP);
UQVB_B49 : OR4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N22, A1 => UQVN_N25, A2 => UQVN_N28, 
	A3 => PS);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => LD);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => CS);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => PS);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => QI4);
UQVB_B54 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N37, A1 => UQVN_N36);
UQVB_B55 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N45, CLK => CLK, CD => CD);
UQVB_B56 : OR4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N38, A1 => UQVN_N39, A2 => UQVN_N35, 
	A3 => PS);
UQVB_B57 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => D4, A1 => LD, A2 => UQVN_N34);
UQVB_B58 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => QI4, A1 => UQVN_N33, A2 => UQVN_N34, 
	A3 => UQVN_N44);
UQVB_B59 : AND9
	PORT MAP (Z0 => UQVN_N39, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => UQVN_N33, A5 => CAI, A6 => EN, 
	A7 => UQVN_N34, A8 => UP);
UQVB_B60 : AND9
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N65, A4 => UQVN_N33, A5 => CAI, A6 => EN, 
	A7 => UQVN_N34, A8 => DNUP);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => QI5);
UQVB_B62 : LXOR2
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N32, A1 => UQVN_N41);
UQVB_B63 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N46, CLK => CLK, CD => CD);
UQVB_B64 : OR4
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N42, A1 => UQVN_N43, A2 => UQVN_N40, 
	A3 => PS);
UQVB_B65 : AND3
	PORT MAP (Z0 => UQVN_N42, A0 => D5, A1 => LD, A2 => UQVN_N34);
UQVB_B66 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => QI5, A1 => UQVN_N33, A2 => UQVN_N34, 
	A3 => UQVN_N44);
UQVB_B67 : AND10
	PORT MAP (Z0 => UQVN_N43, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => UQVN_N33, A6 => CAI, 
	A7 => EN, A8 => UQVN_N34, A9 => UP);
UQVB_B68 : AND10
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N65, A4 => UQVN_N66, A5 => UQVN_N33, A6 => CAI, 
	A7 => EN, A8 => UQVN_N34, A9 => DNUP);
UQVB_B69 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => LD);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => CS);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => PS);
UQVB_B72 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => D6, A1 => LD, A2 => UQVN_N48);
UQVB_B73 : OR4
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N51, A1 => UQVN_N50, A2 => UQVN_N49, 
	A3 => PS);
UQVB_B74 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N60, CLK => CLK, CD => CD);
UQVB_B75 : LXOR2
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N52, A1 => UQVN_N53);
UQVB_B76 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => QI6);
UQVB_B77 : AND4
	PORT MAP (Z0 => UQVN_N52, A0 => QI6, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => UQVN_N54);
UQVB_B78 : AND11
	PORT MAP (Z0 => UQVN_N50, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => UQVN_N47, 
	A7 => CAI, A8 => EN, A9 => UQVN_N48, A10 => UP);
UQVB_B79 : AND11
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N65, A4 => UQVN_N66, A5 => UQVN_N67, A6 => UQVN_N47, 
	A7 => CAI, A8 => EN, A9 => UQVN_N48, A10 => DNUP);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => QI7);
UQVB_B81 : LXOR2
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N58, A1 => UQVN_N57);
UQVB_B82 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N61, CLK => CLK, CD => CD);
UQVB_B83 : OR4
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N59, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => PS);
UQVB_B84 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => D7, A1 => LD, A2 => UQVN_N48);
UQVB_B85 : AND4
	PORT MAP (Z0 => UQVN_N58, A0 => QI7, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => UQVN_N54);
UQVB_B86 : AND12
	PORT MAP (Z0 => UQVN_N56, A0 => QI0, A1 => QI1, A2 => QI2, 
	A3 => QI3, A4 => QI4, A5 => QI5, A6 => QI6, 
	A7 => UQVN_N47, A8 => CAI, A9 => EN, A10 => UQVN_N48, 
	A11 => UP);
UQVB_B87 : AND12
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N65, A4 => UQVN_N66, A5 => UQVN_N67, A6 => UQVN_N68, 
	A7 => UQVN_N47, A8 => CAI, A9 => EN, A10 => UQVN_N48, 
	A11 => DNUP);
END lattice_arch;
-- VHDL netlist for CDD14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CDD14;


ARCHITECTURE lattice_arch OF CDD14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, HOLD0, HOLD1,
	 HOLD2, HOLD3, LOAD0, LOAD1,
	 LOAD2, LOAD3, QI0, QI1,
	 QI2, QI3, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N23, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B2 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N26, A1 => QI2, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B3 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N25, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B5 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B6 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N14);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B8 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N14);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B12 : OR4
	PORT MAP (Z0 => UQVN_N17, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => HOLD0, A1 => UQVN_N8);
UQVB_B18 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD1, A1 => UQVN_N18);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD2, A1 => UQVN_N11);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD3, A1 => UQVN_N17);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI3);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI2);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI1);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI0);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => LD);
UQVB_B26 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B27 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B28 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B29 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B30 : AND2
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N26, A1 => UQVN_N14, A2 => EN);
UQVB_B32 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B33 : AND2
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD);
UQVB_B34 : AND2
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B36 : AND5
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B37 : AND2
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD);
UQVB_B38 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => LOAD2, A1 => UQVN_N16, A2 => UQVN_N19, 
	A3 => UQVN_N15);
UQVB_B39 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N14);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => QI0, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B41 : OR4
	PORT MAP (Z0 => UQVN_N8, A0 => LOAD0, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N22);
UQVB_B42 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N14);
END lattice_arch;
-- VHDL netlist for CDD18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD18 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END CDD18;


ARCHITECTURE lattice_arch OF CDD18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, HOLD0, HOLD1,
	 HOLD2, HOLD3, HOLD4, HOLD5,
	 HOLD6, HOLD7, LOAD0, LOAD1,
	 LOAD2, LOAD3, QI0, QI1,
	 QI2, QI3, QI4, QI5,
	 QI6, QI7, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N51, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B2 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N54, A1 => QI2, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B3 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N53, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B5 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B6 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N14);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B8 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N14);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N53, A1 => UQVN_N52, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B12 : OR4
	PORT MAP (Z0 => UQVN_N17, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => HOLD0, A1 => UQVN_N8);
UQVB_B22 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD1, A1 => UQVN_N18);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD2, A1 => UQVN_N11);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD3, A1 => UQVN_N17);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI3);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => QI2);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => QI1);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI0);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => LD);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B31 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B32 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B33 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B34 : AND2
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N54, A1 => UQVN_N14, A2 => EN);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N53, A1 => UQVN_N52, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B37 : AND2
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD);
UQVB_B38 : AND2
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD);
UQVB_B39 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => UQVN_N52, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B40 : AND5
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N52, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => EN);
UQVB_B41 : AND2
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD);
UQVB_B42 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => LOAD2, A1 => UQVN_N16, A2 => UQVN_N19, 
	A3 => UQVN_N15);
UQVB_B43 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N14);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => QI0, A2 => UQVN_N14, 
	A3 => EN);
UQVB_B45 : OR4
	PORT MAP (Z0 => UQVN_N8, A0 => LOAD0, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N22);
UQVB_B46 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N14);
UQVB_B47 : AND9
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N58, A1 => QI6, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N23, A8 => EN);
UQVB_B48 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N23, A4 => EN);
UQVB_B49 : AND5
	PORT MAP (Z0 => UQVN_N25, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N23, A4 => EN);
UQVB_B50 : OR5
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N31, A1 => UQVN_N32, A2 => UQVN_N33, 
	A3 => UQVN_N24, A4 => UQVN_N25);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => QI7, A1 => QI5, A2 => UQVN_N23, 
	A3 => EN);
UQVB_B52 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => QI5, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N53, A4 => UQVN_N52, A5 => UQVN_N51, A6 => UQVN_N23, 
	A7 => EN);
UQVB_B53 : AND9
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => UQVN_N57, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N23, A8 => EN);
UQVB_B54 : OR5
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N28, A2 => UQVN_N36, 
	A3 => UQVN_N27, A4 => UQVN_N26);
UQVB_B55 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B56 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => HOLD4, A1 => UQVN_N29);
UQVB_B57 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B58 : LXOR2
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD5, A1 => UQVN_N35);
UQVB_B59 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI5);
UQVB_B60 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI4);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => LD);
UQVB_B62 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => D4, A1 => LD);
UQVB_B63 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => D5, A1 => LD);
UQVB_B64 : AND2
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N23);
UQVB_B65 : AND2
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N23);
UQVB_B66 : AND7
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N58, A1 => UQVN_N54, A2 => UQVN_N53, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => UQVN_N23, A6 => EN);
UQVB_B67 : AND8
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N57, A1 => UQVN_N56, A2 => UQVN_N54, 
	A3 => UQVN_N53, A4 => UQVN_N52, A5 => UQVN_N51, A6 => UQVN_N23, 
	A7 => EN);
UQVB_B68 : AND9
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N47, A8 => EN);
UQVB_B69 : AND9
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N57, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N47, A8 => EN);
UQVB_B70 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => QI7, A1 => QI6, A2 => UQVN_N47, 
	A3 => EN);
UQVB_B71 : AND4
	PORT MAP (Z0 => UQVN_N39, A0 => QI7, A1 => QI6, A2 => UQVN_N47, 
	A3 => EN);
UQVB_B72 : AND4
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI5, A2 => UQVN_N47, 
	A3 => EN);
UQVB_B73 : AND9
	PORT MAP (Z0 => UQVN_N43, A0 => QI6, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N47, A8 => EN);
UQVB_B74 : OR4
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N50, A1 => UQVN_N42, A2 => UQVN_N43, 
	A3 => UQVN_N38);
UQVB_B75 : OR4
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N48, A1 => UQVN_N41, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B76 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => HOLD6, A1 => UQVN_N44);
UQVB_B77 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N45, CLK => CLK, CD => CD);
UQVB_B78 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N46, CLK => CLK, CD => CD);
UQVB_B79 : LXOR2
	PORT MAP (Z0 => UQVN_N46, A0 => HOLD7, A1 => UQVN_N49);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => QI7);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => QI6);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => LD);
UQVB_B83 : AND2
	PORT MAP (Z0 => UQVN_N50, A0 => D6, A1 => LD);
UQVB_B84 : AND2
	PORT MAP (Z0 => UQVN_N48, A0 => D7, A1 => LD);
UQVB_B85 : AND2
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N47);
UQVB_B86 : AND2
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N47);
END lattice_arch;
-- VHDL netlist for CDD24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD24 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CDD24;


ARCHITECTURE lattice_arch OF CDD24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, HOLD0,
	 HOLD1, HOLD2, HOLD3, LOAD0,
	 LOAD1, LOAD2, LOAD3, QI0,
	 QI1, QI2, QI3, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => UQVN_N19, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B4 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B5 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N8);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N27, A1 => UQVN_N15, A2 => EN, 
	A3 => UQVN_N8);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI0, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B9 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B10 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N8);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N24, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N27, A1 => QI2, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B13 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N26, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B15 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B16 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N8);
UQVB_B17 : AND6
	PORT MAP (Z0 => UQVN_N17, A0 => QI3, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B18 : AND6
	PORT MAP (Z0 => UQVN_N20, A0 => QI2, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B19 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B20 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B21 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N8);
UQVB_B22 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B23 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B24 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD0, A1 => UQVN_N9);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD1, A1 => UQVN_N19);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD2, A1 => UQVN_N12);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD3, A1 => UQVN_N18);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI0);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => LD);
UQVB_B38 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N10, CLK => CLK);
UQVB_B39 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N11, CLK => CLK);
UQVB_B40 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N13, CLK => CLK);
UQVB_B41 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N14, CLK => CLK);
UQVB_B42 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => LOAD2, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => UQVN_N16);
UQVB_B43 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => LOAD0, A1 => UQVN_N22, A2 => UQVN_N21, 
	A3 => UQVN_N23);
END lattice_arch;
-- VHDL netlist for CDD28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD28 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END CDD28;


ARCHITECTURE lattice_arch OF CDD28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, HOLD0, HOLD1, HOLD2,
	 HOLD3, HOLD4, HOLD5, HOLD6,
	 HOLD7, LOAD0, LOAD1, LOAD2,
	 LOAD3, QI0, QI1, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => UQVN_N19, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B4 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B5 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N8);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N57, A1 => UQVN_N15, A2 => EN, 
	A3 => UQVN_N8);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N56, A1 => UQVN_N55, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI0, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B9 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B10 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N8);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N54, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N57, A1 => QI2, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B13 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N56, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B15 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B16 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N8);
UQVB_B17 : AND6
	PORT MAP (Z0 => UQVN_N17, A0 => QI3, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B18 : AND6
	PORT MAP (Z0 => UQVN_N20, A0 => QI2, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B19 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B20 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B21 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N8);
UQVB_B22 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N56, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => UQVN_N8);
UQVB_B23 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B24 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => UQVN_N8);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD0, A1 => UQVN_N9);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD1, A1 => UQVN_N19);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD2, A1 => UQVN_N12);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD3, A1 => UQVN_N18);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => QI3);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI2);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI1);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI0);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => LD);
UQVB_B42 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N10, CLK => CLK);
UQVB_B43 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N11, CLK => CLK);
UQVB_B44 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N13, CLK => CLK);
UQVB_B45 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N14, CLK => CLK);
UQVB_B46 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => LOAD2, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => UQVN_N16);
UQVB_B47 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => LOAD0, A1 => UQVN_N22, A2 => UQVN_N21, 
	A3 => UQVN_N23);
UQVB_B48 : OR5
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N33, A1 => UQVN_N34, A2 => UQVN_N35, 
	A3 => UQVN_N25, A4 => UQVN_N26);
UQVB_B49 : OR5
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N39, A1 => UQVN_N29, A2 => UQVN_N38, 
	A3 => UQVN_N28, A4 => UQVN_N27);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => CS);
UQVB_B51 : AND3
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N24, A2 => UQVN_N30);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => D4, A1 => LD, A2 => UQVN_N30);
UQVB_B53 : AND8
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N61, A1 => UQVN_N57, A2 => UQVN_N56, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => UQVN_N24, A6 => EN, 
	A7 => UQVN_N30);
UQVB_B54 : AND9
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N60, A1 => UQVN_N59, A2 => UQVN_N57, 
	A3 => UQVN_N56, A4 => UQVN_N55, A5 => UQVN_N54, A6 => UQVN_N24, 
	A7 => EN, A8 => UQVN_N30);
UQVB_B55 : AND6
	PORT MAP (Z0 => UQVN_N25, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N24, A4 => EN, A5 => UQVN_N30);
UQVB_B56 : AND6
	PORT MAP (Z0 => UQVN_N26, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N24, A4 => EN, A5 => UQVN_N30);
UQVB_B57 : AND3
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N24, A2 => UQVN_N30);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => D5, A1 => LD, A2 => UQVN_N30);
UQVB_B59 : AND9
	PORT MAP (Z0 => UQVN_N29, A0 => QI5, A1 => UQVN_N58, A2 => UQVN_N57, 
	A3 => UQVN_N56, A4 => UQVN_N55, A5 => UQVN_N54, A6 => UQVN_N24, 
	A7 => EN, A8 => UQVN_N30);
UQVB_B60 : AND10
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N61, A1 => QI6, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N24, A8 => EN, A9 => UQVN_N30);
UQVB_B61 : AND10
	PORT MAP (Z0 => UQVN_N28, A0 => QI7, A1 => UQVN_N60, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N24, A8 => EN, A9 => UQVN_N30);
UQVB_B62 : AND5
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => QI5, A2 => UQVN_N24, 
	A3 => EN, A4 => UQVN_N30);
UQVB_B63 : FD11
	PORT MAP (Q0 => QI4, D0 => UQVN_N32, CLK => CLK);
UQVB_B64 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => HOLD4, A1 => UQVN_N31);
UQVB_B65 : FD11
	PORT MAP (Q0 => QI5, D0 => UQVN_N36, CLK => CLK);
UQVB_B66 : LXOR2
	PORT MAP (Z0 => UQVN_N36, A0 => HOLD5, A1 => UQVN_N37);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => QI5);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => QI4);
UQVB_B69 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => LD);
UQVB_B70 : OR4
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N53, A1 => UQVN_N44, A2 => UQVN_N45, 
	A3 => UQVN_N40);
UQVB_B71 : OR4
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N51, A1 => UQVN_N43, A2 => UQVN_N41, 
	A3 => UQVN_N42);
UQVB_B72 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => CS);
UQVB_B73 : AND3
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N50, A2 => UQVN_N46);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N53, A0 => D6, A1 => LD, A2 => UQVN_N46);
UQVB_B75 : AND10
	PORT MAP (Z0 => UQVN_N44, A0 => QI7, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N50, A8 => EN, A9 => UQVN_N46);
UQVB_B76 : AND10
	PORT MAP (Z0 => UQVN_N45, A0 => QI6, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N50, A8 => EN, A9 => UQVN_N46);
UQVB_B77 : AND5
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI6, A2 => UQVN_N50, 
	A3 => EN, A4 => UQVN_N46);
UQVB_B78 : AND3
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N50, A2 => UQVN_N46);
UQVB_B79 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => D7, A1 => LD, A2 => UQVN_N46);
UQVB_B80 : AND10
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N60, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N50, A8 => EN, A9 => UQVN_N46);
UQVB_B81 : AND5
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => QI6, A2 => UQVN_N50, 
	A3 => EN, A4 => UQVN_N46);
UQVB_B82 : AND5
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => QI5, A2 => UQVN_N50, 
	A3 => EN, A4 => UQVN_N46);
UQVB_B83 : LXOR2
	PORT MAP (Z0 => UQVN_N48, A0 => HOLD6, A1 => UQVN_N47);
UQVB_B84 : FD11
	PORT MAP (Q0 => QI6, D0 => UQVN_N48, CLK => CLK);
UQVB_B85 : FD11
	PORT MAP (Q0 => QI7, D0 => UQVN_N49, CLK => CLK);
UQVB_B86 : LXOR2
	PORT MAP (Z0 => UQVN_N49, A0 => HOLD7, A1 => UQVN_N52);
UQVB_B87 : INV
	PORT MAP (ZN0 => UQVN_N61, A0 => QI7);
UQVB_B88 : INV
	PORT MAP (ZN0 => UQVN_N60, A0 => QI6);
UQVB_B89 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => LD);
END lattice_arch;
-- VHDL netlist for CDD34
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDD34;


ARCHITECTURE lattice_arch OF CDD34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, HOLD0, HOLD1,
	 HOLD2, HOLD3, LOAD0, LOAD1,
	 LOAD2, LOAD3, QI0, QI1,
	 QI2, QI3, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N14);
UQVB_B3 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N14);
UQVB_B4 : OR4
	PORT MAP (Z0 => UQVN_N17, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N26, A1 => UQVN_N14, A2 => CAI, 
	A3 => EN);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => QI0, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N23, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N26, A1 => QI2, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N25, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B13 : AND6
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B16 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B17 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B18 : AND6
	PORT MAP (Z0 => CAO, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N23, A4 => CAI, A5 => EN);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => HOLD0, A1 => UQVN_N8);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD1, A1 => UQVN_N18);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD2, A1 => UQVN_N11);
UQVB_B26 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD3, A1 => UQVN_N17);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI3);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI2);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI1);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI0);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => LD);
UQVB_B32 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B33 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B34 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B35 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B36 : AND2
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD);
UQVB_B37 : AND2
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD);
UQVB_B38 : AND2
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD);
UQVB_B39 : AND2
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD);
UQVB_B40 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => LOAD2, A1 => UQVN_N16, A2 => UQVN_N19, 
	A3 => UQVN_N15);
UQVB_B41 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N14);
UQVB_B42 : OR4
	PORT MAP (Z0 => UQVN_N8, A0 => LOAD0, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N22);
UQVB_B43 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N14);
END lattice_arch;
-- VHDL netlist for CDD38
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDD38;


ARCHITECTURE lattice_arch OF CDD38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, HOLD0, HOLD1,
	 HOLD2, HOLD3, HOLD4, HOLD5,
	 HOLD6, HOLD7, LOAD0, LOAD1,
	 LOAD2, LOAD3, QI0, QI1,
	 QI2, QI3, QI4, QI5,
	 QI6, QI7, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N14);
UQVB_B3 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N14);
UQVB_B4 : OR4
	PORT MAP (Z0 => UQVN_N17, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N54, A1 => UQVN_N14, A2 => CAI, 
	A3 => EN);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N53, A1 => UQVN_N52, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => QI0, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N51, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N54, A1 => QI2, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N53, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => UQVN_N52, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B13 : AND6
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N52, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N53, A1 => UQVN_N52, A2 => UQVN_N51, 
	A3 => UQVN_N14, A4 => CAI, A5 => EN);
UQVB_B16 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B17 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N14, 
	A3 => CAI, A4 => EN);
UQVB_B18 : AND10
	PORT MAP (Z0 => CAO, A0 => UQVN_N58, A1 => UQVN_N57, A2 => UQVN_N56, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => UQVN_N53, A6 => UQVN_N52, 
	A7 => UQVN_N51, A8 => CAI, A9 => EN);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B27 : LXOR2
	PORT MAP (Z0 => UQVN_N9, A0 => HOLD0, A1 => UQVN_N8);
UQVB_B28 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD1, A1 => UQVN_N18);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD2, A1 => UQVN_N11);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD3, A1 => UQVN_N17);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI3);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => QI2);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => QI1);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI0);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => LD);
UQVB_B36 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B37 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B38 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N12, CLK => CLK, CD => CD);
UQVB_B39 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B40 : AND2
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD);
UQVB_B41 : AND2
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD);
UQVB_B42 : AND2
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD);
UQVB_B43 : AND2
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD);
UQVB_B44 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => LOAD2, A1 => UQVN_N16, A2 => UQVN_N19, 
	A3 => UQVN_N15);
UQVB_B45 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N14);
UQVB_B46 : OR4
	PORT MAP (Z0 => UQVN_N8, A0 => LOAD0, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N22);
UQVB_B47 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N14);
UQVB_B48 : OR5
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N31, A1 => UQVN_N32, A2 => UQVN_N33, 
	A3 => UQVN_N24, A4 => UQVN_N25);
UQVB_B49 : OR5
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N28, A2 => UQVN_N36, 
	A3 => UQVN_N27, A4 => UQVN_N26);
UQVB_B50 : AND8
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N58, A1 => UQVN_N54, A2 => UQVN_N53, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => UQVN_N23, A6 => EN, 
	A7 => CAI);
UQVB_B51 : AND9
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N57, A1 => UQVN_N56, A2 => UQVN_N54, 
	A3 => UQVN_N53, A4 => UQVN_N52, A5 => UQVN_N51, A6 => UQVN_N23, 
	A7 => EN, A8 => CAI);
UQVB_B52 : AND6
	PORT MAP (Z0 => UQVN_N24, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N23, A4 => EN, A5 => CAI);
UQVB_B53 : AND6
	PORT MAP (Z0 => UQVN_N25, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N23, A4 => EN, A5 => CAI);
UQVB_B54 : AND9
	PORT MAP (Z0 => UQVN_N28, A0 => QI5, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N53, A4 => UQVN_N52, A5 => UQVN_N51, A6 => UQVN_N23, 
	A7 => EN, A8 => CAI);
UQVB_B55 : AND10
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N58, A1 => QI6, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N23, A8 => EN, A9 => CAI);
UQVB_B56 : AND10
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => UQVN_N57, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N23, A8 => EN, A9 => CAI);
UQVB_B57 : AND5
	PORT MAP (Z0 => UQVN_N26, A0 => QI7, A1 => QI5, A2 => UQVN_N23, 
	A3 => EN, A4 => CAI);
UQVB_B58 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => HOLD4, A1 => UQVN_N29);
UQVB_B60 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B61 : LXOR2
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD5, A1 => UQVN_N35);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI5);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI4);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => LD);
UQVB_B65 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => D4, A1 => LD);
UQVB_B66 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => D5, A1 => LD);
UQVB_B67 : AND2
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N23);
UQVB_B68 : AND2
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N23);
UQVB_B69 : OR4
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N50, A1 => UQVN_N42, A2 => UQVN_N43, 
	A3 => UQVN_N38);
UQVB_B70 : OR4
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N48, A1 => UQVN_N41, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B71 : AND10
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N47, A8 => EN, A9 => CAI);
UQVB_B72 : AND10
	PORT MAP (Z0 => UQVN_N43, A0 => QI6, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N47, A8 => EN, A9 => CAI);
UQVB_B73 : AND5
	PORT MAP (Z0 => UQVN_N38, A0 => QI7, A1 => QI6, A2 => UQVN_N47, 
	A3 => EN, A4 => CAI);
UQVB_B74 : AND10
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N57, A1 => UQVN_N56, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => UQVN_N53, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => UQVN_N47, A8 => EN, A9 => CAI);
UQVB_B75 : AND5
	PORT MAP (Z0 => UQVN_N39, A0 => QI7, A1 => QI6, A2 => UQVN_N47, 
	A3 => EN, A4 => CAI);
UQVB_B76 : AND5
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI5, A2 => UQVN_N47, 
	A3 => EN, A4 => CAI);
UQVB_B77 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => HOLD6, A1 => UQVN_N44);
UQVB_B78 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N45, CLK => CLK, CD => CD);
UQVB_B79 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N46, CLK => CLK, CD => CD);
UQVB_B80 : LXOR2
	PORT MAP (Z0 => UQVN_N46, A0 => HOLD7, A1 => UQVN_N49);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => QI7);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => QI6);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => LD);
UQVB_B84 : AND2
	PORT MAP (Z0 => UQVN_N50, A0 => D6, A1 => LD);
UQVB_B85 : AND2
	PORT MAP (Z0 => UQVN_N48, A0 => D7, A1 => LD);
UQVB_B86 : AND2
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N47);
UQVB_B87 : AND2
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N47);
END lattice_arch;
-- VHDL netlist for CDD44
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDD44;


ARCHITECTURE lattice_arch OF CDD44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, HOLD0,
	 HOLD1, HOLD2, HOLD3, LOAD0,
	 LOAD1, LOAD2, LOAD3, QI0,
	 QI1, QI2, QI3, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => UQVN_N19, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B3 : AND6
	PORT MAP (Z0 => CAO, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N25, 
	A3 => UQVN_N24, A4 => EN, A5 => CAI);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B5 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B6 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N8);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N27, A1 => UQVN_N15, A2 => EN, 
	A3 => CAI, A4 => UQVN_N8);
UQVB_B8 : AND6
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI0, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B10 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B11 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N8);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N24, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B13 : AND7
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N27, A1 => QI2, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B14 : AND7
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N26, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B16 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B17 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N8);
UQVB_B18 : AND7
	PORT MAP (Z0 => UQVN_N17, A0 => QI3, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B19 : AND7
	PORT MAP (Z0 => UQVN_N20, A0 => QI2, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B20 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B21 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B22 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N8);
UQVB_B23 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B24 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B25 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD0, A1 => UQVN_N9);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD1, A1 => UQVN_N19);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD2, A1 => UQVN_N12);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD3, A1 => UQVN_N18);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI0);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => LD);
UQVB_B39 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N10, CLK => CLK);
UQVB_B40 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N11, CLK => CLK);
UQVB_B41 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N13, CLK => CLK);
UQVB_B42 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N14, CLK => CLK);
UQVB_B43 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => LOAD2, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => UQVN_N16);
UQVB_B44 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => LOAD0, A1 => UQVN_N22, A2 => UQVN_N21, 
	A3 => UQVN_N23);
END lattice_arch;
-- VHDL netlist for CDD48
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDD48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDD48;


ARCHITECTURE lattice_arch OF CDD48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, HOLD0, HOLD1, HOLD2,
	 HOLD3, HOLD4, HOLD5, HOLD6,
	 HOLD7, LOAD0, LOAD1, LOAD2,
	 LOAD3, QI0, QI1, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => UQVN_N19, A0 => LOAD1, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N18, A0 => LOAD3, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N7);
UQVB_B3 : AND10
	PORT MAP (Z0 => CAO, A0 => UQVN_N61, A1 => UQVN_N60, A2 => UQVN_N59, 
	A3 => UQVN_N58, A4 => UQVN_N57, A5 => UQVN_N56, A6 => UQVN_N55, 
	A7 => UQVN_N54, A8 => EN, A9 => CAI);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B5 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B6 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N8);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N57, A1 => UQVN_N15, A2 => EN, 
	A3 => CAI, A4 => UQVN_N8);
UQVB_B8 : AND6
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N56, A1 => UQVN_N55, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI0, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B10 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B11 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N8);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => QI1, A1 => UQVN_N54, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B13 : AND7
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N57, A1 => QI2, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B14 : AND7
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => UQVN_N56, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B16 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B17 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N8);
UQVB_B18 : AND7
	PORT MAP (Z0 => UQVN_N17, A0 => QI3, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B19 : AND7
	PORT MAP (Z0 => UQVN_N20, A0 => QI2, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B20 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B21 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N15, A2 => UQVN_N8);
UQVB_B22 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N8);
UQVB_B23 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N56, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => UQVN_N15, A4 => EN, A5 => CAI, A6 => UQVN_N8);
UQVB_B24 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B25 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N15, 
	A3 => EN, A4 => CAI, A5 => UQVN_N8);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD0, A1 => UQVN_N9);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD1, A1 => UQVN_N19);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD2, A1 => UQVN_N12);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD3, A1 => UQVN_N18);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => QI3);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI2);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI1);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI0);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => LD);
UQVB_B43 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N10, CLK => CLK);
UQVB_B44 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N11, CLK => CLK);
UQVB_B45 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N13, CLK => CLK);
UQVB_B46 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N14, CLK => CLK);
UQVB_B47 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => LOAD2, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => UQVN_N16);
UQVB_B48 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => LOAD0, A1 => UQVN_N22, A2 => UQVN_N21, 
	A3 => UQVN_N23);
UQVB_B49 : OR5
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N33, A1 => UQVN_N34, A2 => UQVN_N35, 
	A3 => UQVN_N25, A4 => UQVN_N26);
UQVB_B50 : OR5
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N39, A1 => UQVN_N29, A2 => UQVN_N38, 
	A3 => UQVN_N28, A4 => UQVN_N27);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => CS);
UQVB_B52 : AND3
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N24, A2 => UQVN_N30);
UQVB_B53 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => D4, A1 => LD, A2 => UQVN_N30);
UQVB_B54 : AND9
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N61, A1 => UQVN_N57, A2 => UQVN_N56, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => UQVN_N24, A6 => EN, 
	A7 => CAI, A8 => UQVN_N30);
UQVB_B55 : AND10
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N60, A1 => UQVN_N59, A2 => UQVN_N57, 
	A3 => UQVN_N56, A4 => UQVN_N55, A5 => UQVN_N54, A6 => UQVN_N24, 
	A7 => EN, A8 => CAI, A9 => UQVN_N30);
UQVB_B56 : AND7
	PORT MAP (Z0 => UQVN_N25, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N24, A4 => EN, A5 => CAI, A6 => UQVN_N30);
UQVB_B57 : AND7
	PORT MAP (Z0 => UQVN_N26, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N24, A4 => EN, A5 => CAI, A6 => UQVN_N30);
UQVB_B58 : AND3
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N24, A2 => UQVN_N30);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => D5, A1 => LD, A2 => UQVN_N30);
UQVB_B60 : AND10
	PORT MAP (Z0 => UQVN_N29, A0 => QI5, A1 => UQVN_N58, A2 => UQVN_N57, 
	A3 => UQVN_N56, A4 => UQVN_N55, A5 => UQVN_N54, A6 => UQVN_N24, 
	A7 => EN, A8 => CAI, A9 => UQVN_N30);
UQVB_B61 : AND11
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N61, A1 => QI6, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N24, A8 => EN, A9 => CAI, A10 => UQVN_N30);
UQVB_B62 : AND11
	PORT MAP (Z0 => UQVN_N28, A0 => QI7, A1 => UQVN_N60, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N24, A8 => EN, A9 => CAI, A10 => UQVN_N30);
UQVB_B63 : AND6
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => QI5, A2 => UQVN_N24, 
	A3 => EN, A4 => CAI, A5 => UQVN_N30);
UQVB_B64 : FD11
	PORT MAP (Q0 => QI4, D0 => UQVN_N32, CLK => CLK);
UQVB_B65 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => HOLD4, A1 => UQVN_N31);
UQVB_B66 : FD11
	PORT MAP (Q0 => QI5, D0 => UQVN_N36, CLK => CLK);
UQVB_B67 : LXOR2
	PORT MAP (Z0 => UQVN_N36, A0 => HOLD5, A1 => UQVN_N37);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => QI5);
UQVB_B69 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => QI4);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => LD);
UQVB_B71 : OR4
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N53, A1 => UQVN_N44, A2 => UQVN_N45, 
	A3 => UQVN_N40);
UQVB_B72 : OR4
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N51, A1 => UQVN_N43, A2 => UQVN_N41, 
	A3 => UQVN_N42);
UQVB_B73 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => CS);
UQVB_B74 : AND3
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N50, A2 => UQVN_N46);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N53, A0 => D6, A1 => LD, A2 => UQVN_N46);
UQVB_B76 : AND11
	PORT MAP (Z0 => UQVN_N44, A0 => QI7, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N50, A8 => EN, A9 => CAI, A10 => UQVN_N46);
UQVB_B77 : AND11
	PORT MAP (Z0 => UQVN_N45, A0 => QI6, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N50, A8 => EN, A9 => CAI, A10 => UQVN_N46);
UQVB_B78 : AND6
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI6, A2 => UQVN_N50, 
	A3 => EN, A4 => CAI, A5 => UQVN_N46);
UQVB_B79 : AND3
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N50, A2 => UQVN_N46);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => D7, A1 => LD, A2 => UQVN_N46);
UQVB_B81 : AND11
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N60, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N56, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => UQVN_N50, A8 => EN, A9 => CAI, A10 => UQVN_N46);
UQVB_B82 : AND6
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => QI6, A2 => UQVN_N50, 
	A3 => EN, A4 => CAI, A5 => UQVN_N46);
UQVB_B83 : AND6
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => QI5, A2 => UQVN_N50, 
	A3 => EN, A4 => CAI, A5 => UQVN_N46);
UQVB_B84 : LXOR2
	PORT MAP (Z0 => UQVN_N48, A0 => HOLD6, A1 => UQVN_N47);
UQVB_B85 : FD11
	PORT MAP (Q0 => QI6, D0 => UQVN_N48, CLK => CLK);
UQVB_B86 : FD11
	PORT MAP (Q0 => QI7, D0 => UQVN_N49, CLK => CLK);
UQVB_B87 : LXOR2
	PORT MAP (Z0 => UQVN_N49, A0 => HOLD7, A1 => UQVN_N52);
UQVB_B88 : INV
	PORT MAP (ZN0 => UQVN_N61, A0 => QI7);
UQVB_B89 : INV
	PORT MAP (ZN0 => UQVN_N60, A0 => QI6);
UQVB_B90 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => LD);
END lattice_arch;
-- VHDL netlist for CDU14
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CDU14;


ARCHITECTURE lattice_arch OF CDU14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 HOLD0, HOLD1, HOLD2, HOLD3,
	 QI0, QI1, QI2, QI3,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N1, A2 => UQVN_N13, 
	A3 => UQVN_N2);
UQVB_B3 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B4 : OR3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N3, A1 => UQVN_N23, A2 => UQVN_N4);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B6 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => UQVN_N24, A2 => UQVN_N5);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B11 : OR5
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N19, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B16 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD0, A1 => UQVN_N10);
UQVB_B18 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B19 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD1, A1 => UQVN_N22);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => HOLD2, A1 => UQVN_N15);
UQVB_B21 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B22 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N17, CLK => CLK, CD => CD);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD3, A1 => UQVN_N20);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => LD);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => D0, A1 => LD);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N27, A1 => UQVN_N18, A2 => EN);
UQVB_B30 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B31 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD);
UQVB_B32 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N27, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => D2, A1 => LD);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D3, A1 => LD);
UQVB_B35 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N18);
UQVB_B36 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N18);
UQVB_B37 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N18);
UQVB_B38 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N27, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN);
UQVB_B39 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N18);
END lattice_arch;
-- VHDL netlist for CDU18
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU18 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END CDU18;


ARCHITECTURE lattice_arch OF CDU18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, HOLD0, HOLD1,
	 HOLD2, HOLD3, HOLD4, HOLD5,
	 HOLD6, HOLD7, QI0, QI1,
	 QI2, QI3, QI4, QI5,
	 QI6, QI7, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N1, A2 => UQVN_N13, 
	A3 => UQVN_N2);
UQVB_B3 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B4 : OR3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N3, A1 => UQVN_N23, A2 => UQVN_N4);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B6 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => UQVN_N24, A2 => UQVN_N5);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B11 : OR5
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N19, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B20 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD0, A1 => UQVN_N10);
UQVB_B22 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD1, A1 => UQVN_N22);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => HOLD2, A1 => UQVN_N15);
UQVB_B25 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B26 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N17, CLK => CLK, CD => CD);
UQVB_B27 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD3, A1 => UQVN_N20);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => QI3);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => QI2);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI1);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => LD);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => D0, A1 => LD);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N53, A1 => UQVN_N18, A2 => EN);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N52, A1 => UQVN_N51, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B35 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N53, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => D2, A1 => LD);
UQVB_B38 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D3, A1 => LD);
UQVB_B39 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N18);
UQVB_B40 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N18);
UQVB_B41 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N18);
UQVB_B42 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N53, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN);
UQVB_B43 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N18);
UQVB_B44 : AND8
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N56, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => QI0, A6 => UQVN_N25, 
	A7 => EN);
UQVB_B45 : AND5
	PORT MAP (Z0 => UQVN_N26, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N25, A4 => EN);
UQVB_B46 : AND5
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N25, A4 => EN);
UQVB_B47 : OR5
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N31, A1 => UQVN_N32, A2 => UQVN_N33, 
	A3 => UQVN_N26, A4 => UQVN_N27);
UQVB_B48 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => QI7, A1 => QI5, A2 => UQVN_N25, 
	A3 => EN);
UQVB_B49 : OR3
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N28);
UQVB_B50 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B51 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => HOLD4, A1 => UQVN_N29);
UQVB_B52 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B53 : LXOR2
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD5, A1 => UQVN_N35);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI5);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => LD);
UQVB_B56 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => D4, A1 => LD);
UQVB_B57 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => D5, A1 => LD);
UQVB_B58 : AND2
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N25);
UQVB_B59 : AND2
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N25);
UQVB_B60 : AND7
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N56, A1 => QI3, A2 => UQVN_N52, 
	A3 => UQVN_N51, A4 => QI0, A5 => UQVN_N25, A6 => EN);
UQVB_B61 : AND8
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N55, A1 => UQVN_N54, A2 => QI3, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => QI0, A6 => UQVN_N25, 
	A7 => EN);
UQVB_B62 : AND9
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N56, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N52, A5 => UQVN_N51, A6 => QI0, 
	A7 => UQVN_N46, A8 => EN);
UQVB_B63 : AND9
	PORT MAP (Z0 => UQVN_N42, A0 => QI6, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N52, A5 => UQVN_N51, A6 => QI0, 
	A7 => UQVN_N46, A8 => EN);
UQVB_B64 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => QI7, A1 => QI6, A2 => UQVN_N46, 
	A3 => EN);
UQVB_B65 : OR3
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N49, A1 => UQVN_N50, A2 => UQVN_N38);
UQVB_B66 : AND4
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI6, A2 => UQVN_N46, 
	A3 => EN);
UQVB_B67 : AND4
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => QI5, A2 => UQVN_N46, 
	A3 => EN);
UQVB_B68 : OR5
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N47, A1 => UQVN_N42, A2 => UQVN_N39, 
	A3 => UQVN_N40, A4 => UQVN_N41);
UQVB_B69 : LXOR2
	PORT MAP (Z0 => UQVN_N44, A0 => HOLD6, A1 => UQVN_N43);
UQVB_B70 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N44, CLK => CLK, CD => CD);
UQVB_B71 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N45, CLK => CLK, CD => CD);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => HOLD7, A1 => UQVN_N48);
UQVB_B73 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI7);
UQVB_B74 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI6);
UQVB_B75 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => LD);
UQVB_B76 : AND2
	PORT MAP (Z0 => UQVN_N49, A0 => D6, A1 => LD);
UQVB_B77 : AND2
	PORT MAP (Z0 => UQVN_N47, A0 => D7, A1 => LD);
UQVB_B78 : AND8
	PORT MAP (Z0 => UQVN_N39, A0 => QI7, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => QI0, A6 => UQVN_N46, 
	A7 => EN);
UQVB_B79 : AND2
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N46);
UQVB_B80 : AND2
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N46);
END lattice_arch;
-- VHDL netlist for CDU24
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU24 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CDU24;


ARCHITECTURE lattice_arch OF CDU24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, HOLD0, HOLD1, HOLD2,
	 HOLD3, QI0, QI1, QI2,
	 QI3, UQVN_N26, UQVN_N27, UQVN_N28 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N13, A1 => UQVN_N1, A2 => UQVN_N14, 
	A3 => UQVN_N2);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N3, A1 => UQVN_N24, A2 => UQVN_N4);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N22, A1 => UQVN_N25, A2 => UQVN_N5);
UQVB_B4 : OR5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N20, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B6 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N28, A1 => UQVN_N19, A2 => EN, 
	A3 => UQVN_N10);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B11 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N28, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B15 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D2, A1 => LD, A2 => UQVN_N10);
UQVB_B17 : AND6
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N28, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => UQVN_N10);
UQVB_B18 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B19 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => D3, A1 => LD, A2 => UQVN_N10);
UQVB_B21 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => UQVN_N10);
UQVB_B22 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B23 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B24 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B29 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N12, CLK => CLK);
UQVB_B30 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD0, A1 => UQVN_N11);
UQVB_B31 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N15, CLK => CLK);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => HOLD1, A1 => UQVN_N23);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD2, A1 => UQVN_N16);
UQVB_B34 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N17, CLK => CLK);
UQVB_B35 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N18, CLK => CLK);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N18, A0 => HOLD3, A1 => UQVN_N21);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => QI3);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI2);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI1);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => LD);
END lattice_arch;
-- VHDL netlist for CDU28
-- Date: 15.5.95 13.45.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU28 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END CDU28;


ARCHITECTURE lattice_arch OF CDU28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, HOLD0, HOLD1, HOLD2,
	 HOLD3, HOLD4, HOLD5, HOLD6,
	 HOLD7, QI0, QI1, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N13, A1 => UQVN_N1, A2 => UQVN_N14, 
	A3 => UQVN_N2);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N3, A1 => UQVN_N24, A2 => UQVN_N4);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N22, A1 => UQVN_N25, A2 => UQVN_N5);
UQVB_B4 : OR5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N20, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B6 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N56, A1 => UQVN_N19, A2 => EN, 
	A3 => UQVN_N10);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N55, A1 => UQVN_N54, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B11 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N56, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B15 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D2, A1 => LD, A2 => UQVN_N10);
UQVB_B17 : AND6
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N56, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => UQVN_N10);
UQVB_B18 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B19 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => D3, A1 => LD, A2 => UQVN_N10);
UQVB_B21 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => UQVN_N10);
UQVB_B22 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B23 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B24 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B33 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N12, CLK => CLK);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD0, A1 => UQVN_N11);
UQVB_B35 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N15, CLK => CLK);
UQVB_B36 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => HOLD1, A1 => UQVN_N23);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD2, A1 => UQVN_N16);
UQVB_B38 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N17, CLK => CLK);
UQVB_B39 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N18, CLK => CLK);
UQVB_B40 : LXOR2
	PORT MAP (Z0 => UQVN_N18, A0 => HOLD3, A1 => UQVN_N21);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI3);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI2);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI1);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => LD);
UQVB_B45 : OR5
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N33, A1 => UQVN_N34, A2 => UQVN_N35, 
	A3 => UQVN_N27, A4 => UQVN_N28);
UQVB_B46 : OR3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N39, A1 => UQVN_N38, A2 => UQVN_N29);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => CS);
UQVB_B48 : AND3
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N26, A2 => UQVN_N30);
UQVB_B49 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => D4, A1 => LD, A2 => UQVN_N30);
UQVB_B50 : AND8
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N59, A1 => QI3, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => QI0, A5 => UQVN_N26, A6 => EN, 
	A7 => UQVN_N30);
UQVB_B51 : AND9
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N58, A1 => UQVN_N57, A2 => QI3, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => QI0, A6 => UQVN_N26, 
	A7 => EN, A8 => UQVN_N30);
UQVB_B52 : AND6
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N26, A4 => EN, A5 => UQVN_N30);
UQVB_B53 : AND6
	PORT MAP (Z0 => UQVN_N28, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N26, A4 => EN, A5 => UQVN_N30);
UQVB_B54 : AND3
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N26, A2 => UQVN_N30);
UQVB_B55 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => D5, A1 => LD, A2 => UQVN_N30);
UQVB_B56 : AND9
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N59, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => QI0, A6 => UQVN_N26, 
	A7 => EN, A8 => UQVN_N30);
UQVB_B57 : AND5
	PORT MAP (Z0 => UQVN_N29, A0 => QI7, A1 => QI5, A2 => UQVN_N26, 
	A3 => EN, A4 => UQVN_N30);
UQVB_B58 : FD11
	PORT MAP (Q0 => QI4, D0 => UQVN_N32, CLK => CLK);
UQVB_B59 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => HOLD4, A1 => UQVN_N31);
UQVB_B60 : FD11
	PORT MAP (Q0 => QI5, D0 => UQVN_N36, CLK => CLK);
UQVB_B61 : LXOR2
	PORT MAP (Z0 => UQVN_N36, A0 => HOLD5, A1 => UQVN_N37);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => QI5);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => LD);
UQVB_B64 : OR3
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N52, A1 => UQVN_N53, A2 => UQVN_N40);
UQVB_B65 : OR5
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N50, A1 => UQVN_N44, A2 => UQVN_N41, 
	A3 => UQVN_N42, A4 => UQVN_N43);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => CS);
UQVB_B67 : AND3
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N49, A2 => UQVN_N45);
UQVB_B68 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => D6, A1 => LD, A2 => UQVN_N45);
UQVB_B69 : AND10
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N59, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N55, A5 => UQVN_N54, A6 => QI0, 
	A7 => UQVN_N49, A8 => EN, A9 => UQVN_N45);
UQVB_B70 : AND5
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI6, A2 => UQVN_N49, 
	A3 => EN, A4 => UQVN_N45);
UQVB_B71 : AND3
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N49, A2 => UQVN_N45);
UQVB_B72 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => D7, A1 => LD, A2 => UQVN_N45);
UQVB_B73 : AND10
	PORT MAP (Z0 => UQVN_N44, A0 => QI6, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N55, A5 => UQVN_N54, A6 => QI0, 
	A7 => UQVN_N49, A8 => EN, A9 => UQVN_N45);
UQVB_B74 : AND9
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => QI0, A6 => UQVN_N49, 
	A7 => EN, A8 => UQVN_N45);
UQVB_B75 : AND5
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => QI6, A2 => UQVN_N49, 
	A3 => EN, A4 => UQVN_N45);
UQVB_B76 : AND5
	PORT MAP (Z0 => UQVN_N43, A0 => QI7, A1 => QI5, A2 => UQVN_N49, 
	A3 => EN, A4 => UQVN_N45);
UQVB_B77 : LXOR2
	PORT MAP (Z0 => UQVN_N47, A0 => HOLD6, A1 => UQVN_N46);
UQVB_B78 : FD11
	PORT MAP (Q0 => QI6, D0 => UQVN_N47, CLK => CLK);
UQVB_B79 : FD11
	PORT MAP (Q0 => QI7, D0 => UQVN_N48, CLK => CLK);
UQVB_B80 : LXOR2
	PORT MAP (Z0 => UQVN_N48, A0 => HOLD7, A1 => UQVN_N51);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => QI7);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => QI6);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => LD);
END lattice_arch;
-- VHDL netlist for CDU34
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDU34;


ARCHITECTURE lattice_arch OF CDU34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 HOLD0, HOLD1, HOLD2, HOLD3,
	 QI0, QI1, QI2, QI3,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N1, A2 => UQVN_N13, 
	A3 => UQVN_N2);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N3, A1 => UQVN_N23, A2 => UQVN_N4);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => UQVN_N24, A2 => UQVN_N5);
UQVB_B4 : OR5
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N19, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N27, A1 => UQVN_N18, A2 => EN, 
	A3 => CAI);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N27, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N27, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN, A5 => CAI);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN, A5 => CAI);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B16 : AND6
	PORT MAP (Z0 => CAO, A0 => QI3, A1 => UQVN_N26, A2 => UQVN_N25, 
	A3 => QI0, A4 => EN, A5 => CAI);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B21 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B22 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD0, A1 => UQVN_N10);
UQVB_B23 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD1, A1 => UQVN_N22);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => HOLD2, A1 => UQVN_N15);
UQVB_B26 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B27 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N17, CLK => CLK, CD => CD);
UQVB_B28 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD3, A1 => UQVN_N20);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => LD);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => D0, A1 => LD);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD);
UQVB_B35 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => D2, A1 => LD);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D3, A1 => LD);
UQVB_B37 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N18);
UQVB_B38 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N18);
UQVB_B39 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N18);
UQVB_B40 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N18);
END lattice_arch;
-- VHDL netlist for CDU38
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDU38;


ARCHITECTURE lattice_arch OF CDU38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, HOLD0, HOLD1,
	 HOLD2, HOLD3, HOLD4, HOLD5,
	 HOLD6, HOLD7, QI0, QI1,
	 QI2, QI3, QI4, QI5,
	 QI6, QI7, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N1, A2 => UQVN_N13, 
	A3 => UQVN_N2);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N3, A1 => UQVN_N23, A2 => UQVN_N4);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => UQVN_N24, A2 => UQVN_N5);
UQVB_B4 : OR5
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N19, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N53, A1 => UQVN_N18, A2 => EN, 
	A3 => CAI);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N52, A1 => UQVN_N51, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N53, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N53, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN, A5 => CAI);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N18, A4 => EN, A5 => CAI);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N18, 
	A3 => EN, A4 => CAI);
UQVB_B16 : AND10
	PORT MAP (Z0 => CAO, A0 => QI7, A1 => UQVN_N55, A2 => UQVN_N54, 
	A3 => QI4, A4 => QI3, A5 => UQVN_N52, A6 => UQVN_N51, 
	A7 => QI0, A8 => EN, A9 => CAI);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B25 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B26 : LXOR2
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD0, A1 => UQVN_N10);
UQVB_B27 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B28 : LXOR2
	PORT MAP (Z0 => UQVN_N14, A0 => HOLD1, A1 => UQVN_N22);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => UQVN_N16, A0 => HOLD2, A1 => UQVN_N15);
UQVB_B30 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B31 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N17, CLK => CLK, CD => CD);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD3, A1 => UQVN_N20);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => QI3);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => QI2);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => QI1);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => LD);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => D0, A1 => LD);
UQVB_B38 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD);
UQVB_B39 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => D2, A1 => LD);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D3, A1 => LD);
UQVB_B41 : AND2
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N18);
UQVB_B42 : AND2
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N18);
UQVB_B43 : AND2
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N18);
UQVB_B44 : AND2
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N18);
UQVB_B45 : OR5
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N31, A1 => UQVN_N32, A2 => UQVN_N33, 
	A3 => UQVN_N26, A4 => UQVN_N27);
UQVB_B46 : OR3
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N28);
UQVB_B47 : AND8
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N56, A1 => QI3, A2 => UQVN_N52, 
	A3 => UQVN_N51, A4 => QI0, A5 => UQVN_N25, A6 => EN, 
	A7 => CAI);
UQVB_B48 : AND9
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N55, A1 => UQVN_N54, A2 => QI3, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => QI0, A6 => UQVN_N25, 
	A7 => EN, A8 => CAI);
UQVB_B49 : AND6
	PORT MAP (Z0 => UQVN_N26, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N25, A4 => EN, A5 => CAI);
UQVB_B50 : AND6
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N25, A4 => EN, A5 => CAI);
UQVB_B51 : AND9
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N56, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => QI0, A6 => UQVN_N25, 
	A7 => EN, A8 => CAI);
UQVB_B52 : AND5
	PORT MAP (Z0 => UQVN_N28, A0 => QI7, A1 => QI5, A2 => UQVN_N25, 
	A3 => EN, A4 => CAI);
UQVB_B53 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B54 : LXOR2
	PORT MAP (Z0 => UQVN_N30, A0 => HOLD4, A1 => UQVN_N29);
UQVB_B55 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B56 : LXOR2
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD5, A1 => UQVN_N35);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI5);
UQVB_B58 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => LD);
UQVB_B59 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => D4, A1 => LD);
UQVB_B60 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => D5, A1 => LD);
UQVB_B61 : AND2
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N25);
UQVB_B62 : AND2
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N25);
UQVB_B63 : OR3
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N49, A1 => UQVN_N50, A2 => UQVN_N38);
UQVB_B64 : OR5
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N47, A1 => UQVN_N42, A2 => UQVN_N39, 
	A3 => UQVN_N40, A4 => UQVN_N41);
UQVB_B65 : AND10
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N56, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N52, A5 => UQVN_N51, A6 => QI0, 
	A7 => UQVN_N46, A8 => EN, A9 => CAI);
UQVB_B66 : AND5
	PORT MAP (Z0 => UQVN_N38, A0 => QI7, A1 => QI6, A2 => UQVN_N46, 
	A3 => EN, A4 => CAI);
UQVB_B67 : AND10
	PORT MAP (Z0 => UQVN_N42, A0 => QI6, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N52, A5 => UQVN_N51, A6 => QI0, 
	A7 => UQVN_N46, A8 => EN, A9 => CAI);
UQVB_B68 : AND9
	PORT MAP (Z0 => UQVN_N39, A0 => QI7, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N52, A4 => UQVN_N51, A5 => QI0, A6 => UQVN_N46, 
	A7 => EN, A8 => CAI);
UQVB_B69 : AND5
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI6, A2 => UQVN_N46, 
	A3 => EN, A4 => CAI);
UQVB_B70 : AND5
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => QI5, A2 => UQVN_N46, 
	A3 => EN, A4 => CAI);
UQVB_B71 : LXOR2
	PORT MAP (Z0 => UQVN_N44, A0 => HOLD6, A1 => UQVN_N43);
UQVB_B72 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N44, CLK => CLK, CD => CD);
UQVB_B73 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N45, CLK => CLK, CD => CD);
UQVB_B74 : LXOR2
	PORT MAP (Z0 => UQVN_N45, A0 => HOLD7, A1 => UQVN_N48);
UQVB_B75 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI7);
UQVB_B76 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI6);
UQVB_B77 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => LD);
UQVB_B78 : AND2
	PORT MAP (Z0 => UQVN_N49, A0 => D6, A1 => LD);
UQVB_B79 : AND2
	PORT MAP (Z0 => UQVN_N47, A0 => D7, A1 => LD);
UQVB_B80 : AND2
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N46);
UQVB_B81 : AND2
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N46);
END lattice_arch;
-- VHDL netlist for CDU44
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDU44;


ARCHITECTURE lattice_arch OF CDU44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, HOLD0, HOLD1, HOLD2,
	 HOLD3, QI0, QI1, QI2,
	 QI3, UQVN_N26, UQVN_N27, UQVN_N28 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N13, A1 => UQVN_N1, A2 => UQVN_N14, 
	A3 => UQVN_N2);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N3, A1 => UQVN_N24, A2 => UQVN_N4);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N22, A1 => UQVN_N25, A2 => UQVN_N5);
UQVB_B4 : OR5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N20, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B5 : AND6
	PORT MAP (Z0 => CAO, A0 => QI3, A1 => UQVN_N27, A2 => UQVN_N26, 
	A3 => QI0, A4 => EN, A5 => CAI);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B7 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N28, A1 => UQVN_N19, A2 => EN, 
	A3 => CAI, A4 => UQVN_N10);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B11 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B12 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B14 : AND6
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N28, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D2, A1 => LD, A2 => UQVN_N10);
UQVB_B18 : AND7
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N28, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => CAI, A6 => UQVN_N10);
UQVB_B19 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B20 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => D3, A1 => LD, A2 => UQVN_N10);
UQVB_B22 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => CAI, A6 => UQVN_N10);
UQVB_B23 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B24 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B25 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B30 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N12, CLK => CLK);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD0, A1 => UQVN_N11);
UQVB_B32 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N15, CLK => CLK);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => HOLD1, A1 => UQVN_N23);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD2, A1 => UQVN_N16);
UQVB_B35 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N17, CLK => CLK);
UQVB_B36 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N18, CLK => CLK);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N18, A0 => HOLD3, A1 => UQVN_N21);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => QI3);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI2);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI1);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => LD);
END lattice_arch;
-- VHDL netlist for CDU48
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDU48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDU48;


ARCHITECTURE lattice_arch OF CDU48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, HOLD0, HOLD1, HOLD2,
	 HOLD3, HOLD4, HOLD5, HOLD6,
	 HOLD7, QI0, QI1, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N13, A1 => UQVN_N1, A2 => UQVN_N14, 
	A3 => UQVN_N2);
UQVB_B2 : OR3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N3, A1 => UQVN_N24, A2 => UQVN_N4);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N22, A1 => UQVN_N25, A2 => UQVN_N5);
UQVB_B4 : OR5
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N20, A1 => UQVN_N9, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8);
UQVB_B5 : AND10
	PORT MAP (Z0 => CAO, A0 => QI7, A1 => UQVN_N58, A2 => UQVN_N57, 
	A3 => QI4, A4 => QI3, A5 => UQVN_N55, A6 => UQVN_N54, 
	A7 => QI0, A8 => EN, A9 => CAI);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B7 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N56, A1 => UQVN_N19, A2 => EN, 
	A3 => CAI, A4 => UQVN_N10);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N55, A1 => UQVN_N54, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B11 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B12 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B14 : AND6
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N56, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D2, A1 => LD, A2 => UQVN_N10);
UQVB_B18 : AND7
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N56, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => CAI, A6 => UQVN_N10);
UQVB_B19 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B20 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N19, A2 => UQVN_N10);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => D3, A1 => LD, A2 => UQVN_N10);
UQVB_B22 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N19, A4 => EN, A5 => CAI, A6 => UQVN_N10);
UQVB_B23 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B24 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B25 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => QI2, A2 => UQVN_N19, 
	A3 => EN, A4 => CAI, A5 => UQVN_N10);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B34 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N12, CLK => CLK);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD0, A1 => UQVN_N11);
UQVB_B36 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N15, CLK => CLK);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => UQVN_N15, A0 => HOLD1, A1 => UQVN_N23);
UQVB_B38 : LXOR2
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD2, A1 => UQVN_N16);
UQVB_B39 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N17, CLK => CLK);
UQVB_B40 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N18, CLK => CLK);
UQVB_B41 : LXOR2
	PORT MAP (Z0 => UQVN_N18, A0 => HOLD3, A1 => UQVN_N21);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => QI3);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => QI2);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => QI1);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => LD);
UQVB_B46 : OR5
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N33, A1 => UQVN_N34, A2 => UQVN_N35, 
	A3 => UQVN_N27, A4 => UQVN_N28);
UQVB_B47 : OR3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N39, A1 => UQVN_N38, A2 => UQVN_N29);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => CS);
UQVB_B49 : AND3
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N26, A2 => UQVN_N30);
UQVB_B50 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => D4, A1 => LD, A2 => UQVN_N30);
UQVB_B51 : AND9
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N59, A1 => QI3, A2 => UQVN_N55, 
	A3 => UQVN_N54, A4 => QI0, A5 => UQVN_N26, A6 => EN, 
	A7 => CAI, A8 => UQVN_N30);
UQVB_B52 : AND10
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N58, A1 => UQVN_N57, A2 => QI3, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => QI0, A6 => UQVN_N26, 
	A7 => EN, A8 => CAI, A9 => UQVN_N30);
UQVB_B53 : AND7
	PORT MAP (Z0 => UQVN_N27, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N26, A4 => EN, A5 => CAI, A6 => UQVN_N30);
UQVB_B54 : AND7
	PORT MAP (Z0 => UQVN_N28, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N26, A4 => EN, A5 => CAI, A6 => UQVN_N30);
UQVB_B55 : AND3
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N26, A2 => UQVN_N30);
UQVB_B56 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => D5, A1 => LD, A2 => UQVN_N30);
UQVB_B57 : AND10
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N59, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => QI0, A6 => UQVN_N26, 
	A7 => EN, A8 => CAI, A9 => UQVN_N30);
UQVB_B58 : AND6
	PORT MAP (Z0 => UQVN_N29, A0 => QI7, A1 => QI5, A2 => UQVN_N26, 
	A3 => EN, A4 => CAI, A5 => UQVN_N30);
UQVB_B59 : FD11
	PORT MAP (Q0 => QI4, D0 => UQVN_N32, CLK => CLK);
UQVB_B60 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => HOLD4, A1 => UQVN_N31);
UQVB_B61 : FD11
	PORT MAP (Q0 => QI5, D0 => UQVN_N36, CLK => CLK);
UQVB_B62 : LXOR2
	PORT MAP (Z0 => UQVN_N36, A0 => HOLD5, A1 => UQVN_N37);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => QI5);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => LD);
UQVB_B65 : OR3
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N52, A1 => UQVN_N53, A2 => UQVN_N40);
UQVB_B66 : OR5
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N50, A1 => UQVN_N44, A2 => UQVN_N41, 
	A3 => UQVN_N42, A4 => UQVN_N43);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => CS);
UQVB_B68 : AND3
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N49, A2 => UQVN_N45);
UQVB_B69 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => D6, A1 => LD, A2 => UQVN_N45);
UQVB_B70 : AND11
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N59, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N55, A5 => UQVN_N54, A6 => QI0, 
	A7 => UQVN_N49, A8 => EN, A9 => CAI, A10 => UQVN_N45);
UQVB_B71 : AND6
	PORT MAP (Z0 => UQVN_N40, A0 => QI7, A1 => QI6, A2 => UQVN_N49, 
	A3 => EN, A4 => CAI, A5 => UQVN_N45);
UQVB_B72 : AND3
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N49, A2 => UQVN_N45);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => D7, A1 => LD, A2 => UQVN_N45);
UQVB_B74 : AND11
	PORT MAP (Z0 => UQVN_N44, A0 => QI6, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N55, A5 => UQVN_N54, A6 => QI0, 
	A7 => UQVN_N49, A8 => EN, A9 => CAI, A10 => UQVN_N45);
UQVB_B75 : AND10
	PORT MAP (Z0 => UQVN_N41, A0 => QI7, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N55, A4 => UQVN_N54, A5 => QI0, A6 => UQVN_N49, 
	A7 => EN, A8 => CAI, A9 => UQVN_N45);
UQVB_B76 : AND6
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => QI6, A2 => UQVN_N49, 
	A3 => EN, A4 => CAI, A5 => UQVN_N45);
UQVB_B77 : AND6
	PORT MAP (Z0 => UQVN_N43, A0 => QI7, A1 => QI5, A2 => UQVN_N49, 
	A3 => EN, A4 => CAI, A5 => UQVN_N45);
UQVB_B78 : LXOR2
	PORT MAP (Z0 => UQVN_N47, A0 => HOLD6, A1 => UQVN_N46);
UQVB_B79 : FD11
	PORT MAP (Q0 => QI6, D0 => UQVN_N47, CLK => CLK);
UQVB_B80 : FD11
	PORT MAP (Q0 => QI7, D0 => UQVN_N48, CLK => CLK);
UQVB_B81 : LXOR2
	PORT MAP (Z0 => UQVN_N48, A0 => HOLD7, A1 => UQVN_N51);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => QI7);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => QI6);
UQVB_B84 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => LD);
END lattice_arch;
-- VHDL netlist for CDUD4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDUD4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CDUD4;


ARCHITECTURE lattice_arch OF CDUD4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 HOLD0, HOLD1, HOLD2, HOLD3,
	 LOAD0, LOAD1, LOAD2, QI0,
	 QI1, QI2, QI3, UQVN_N33,
	 UQVN_N34, UQVN_N35, UQVN_N36 : std_logic;


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


BEGIN

UQVB_B1 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => QI0, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N4, A0 => LOAD0, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B3 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N11, A2 => UQVN_N10);
UQVB_B4 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => QI1, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B9 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B10 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B11 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B12 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => HOLD0, A1 => UQVN_N4);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N36, A1 => UQVN_N11, A2 => EN, 
	A3 => UQVN_N10);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N35, A1 => UQVN_N34, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B15 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N6, A0 => HOLD1, A1 => UQVN_N15);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => QI1);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => QI0);
UQVB_B19 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N36, A1 => QI0, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N12, A5 => UQVN_N10);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => LD);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B22 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => QI1, A1 => UQVN_N33, A2 => UQVN_N11, 
	A3 => EN, A4 => DNUP, A5 => UQVN_N10);
UQVB_B23 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N36, A1 => QI2, A2 => UQVN_N33, 
	A3 => UQVN_N11, A4 => EN, A5 => DNUP, A6 => UQVN_N10);
UQVB_B24 : AND7
	PORT MAP (Z0 => UQVN_N13, A0 => QI3, A1 => UQVN_N35, A2 => UQVN_N33, 
	A3 => UQVN_N11, A4 => EN, A5 => DNUP, A6 => UQVN_N10);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => DNUP);
UQVB_B26 : OR6
	PORT MAP (Z0 => UQVN_N15, A0 => LOAD1, A1 => UQVN_N7, A2 => UQVN_N8, 
	A3 => UQVN_N9, A4 => UQVN_N13, A5 => UQVN_N14);
UQVB_B27 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N11, A2 => UQVN_N10);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => LD);
UQVB_B29 : AND7
	PORT MAP (Z0 => UQVN_N17, A0 => QI2, A1 => UQVN_N34, A2 => UQVN_N33, 
	A3 => UQVN_N28, A4 => EN, A5 => DNUP, A6 => UQVN_N29);
UQVB_B30 : AND5
	PORT MAP (Z0 => UQVN_N18, A0 => QI3, A1 => QI2, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N29);
UQVB_B31 : OR5
	PORT MAP (Z0 => UQVN_N22, A0 => LOAD2, A1 => UQVN_N24, A2 => UQVN_N16, 
	A3 => UQVN_N17, A4 => UQVN_N18);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => CS);
UQVB_B33 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N28, A2 => UQVN_N29);
UQVB_B34 : AND5
	PORT MAP (Z0 => UQVN_N27, A0 => QI3, A1 => QI2, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N29);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N30, A0 => QI3, A1 => QI1, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N29);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => DNUP);
UQVB_B37 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N29);
UQVB_B38 : AND7
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N36, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N28, A4 => EN, A5 => UQVN_N25, A6 => UQVN_N29);
UQVB_B39 : OR6
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N19, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N26, A4 => UQVN_N27, A5 => UQVN_N30);
UQVB_B40 : AND7
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => UQVN_N34, A2 => UQVN_N33, 
	A3 => UQVN_N28, A4 => EN, A5 => DNUP, A6 => UQVN_N29);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => D3, A1 => LD, A2 => UQVN_N29);
UQVB_B42 : AND7
	PORT MAP (Z0 => UQVN_N20, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N28, A4 => EN, A5 => UQVN_N25, A6 => UQVN_N29);
UQVB_B43 : AND6
	PORT MAP (Z0 => UQVN_N21, A0 => QI3, A1 => QI0, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N25, A5 => UQVN_N29);
UQVB_B44 : AND7
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N35, A1 => UQVN_N34, A2 => UQVN_N33, 
	A3 => UQVN_N28, A4 => EN, A5 => DNUP, A6 => UQVN_N29);
UQVB_B45 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => HOLD3, A1 => UQVN_N31);
UQVB_B46 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => HOLD2, A1 => UQVN_N22);
UQVB_B47 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N32, CLK => CLK, CD => CD);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => QI2);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => QI3);
UQVB_B50 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B51 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N28, A2 => UQVN_N29);
END lattice_arch;
-- VHDL netlist for CDUD4C
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDUD4C IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDUD4C;


ARCHITECTURE lattice_arch OF CDUD4C IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, HOLD0, HOLD1,
	 HOLD2, HOLD3, LOAD0, LOAD1,
	 LOAD2, QI0, QI1, QI2,
	 QI3, UQVN_N35, UQVN_N36, UQVN_N37,
	 UQVN_N38 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N6, A0 => LOAD0, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B2 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N13, A2 => UQVN_N12);
UQVB_B3 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N38, A1 => UQVN_N13, A2 => EN, 
	A3 => CAI, A4 => UQVN_N12);
UQVB_B4 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N12);
UQVB_B5 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => QI0, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N12);
UQVB_B6 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N38, A1 => QI0, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N14, A6 => UQVN_N12);
UQVB_B7 : AND7
	PORT MAP (Z0 => UQVN_N10, A0 => QI1, A1 => UQVN_N35, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => DNUP, A6 => UQVN_N12);
UQVB_B8 : AND8
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N38, A1 => QI2, A2 => UQVN_N35, 
	A3 => UQVN_N13, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N12);
UQVB_B9 : AND8
	PORT MAP (Z0 => UQVN_N15, A0 => QI3, A1 => UQVN_N37, A2 => UQVN_N35, 
	A3 => UQVN_N13, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N12);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI1, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N12);
UQVB_B11 : AND7
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35, A4 => EN, A5 => CAI, A6 => DNUP);
UQVB_B12 : AND7
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => QI0, A4 => EN, A5 => CAI, A6 => UQVN_N14);
UQVB_B13 : OR2
	PORT MAP (Z0 => CAO, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B18 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N12);
UQVB_B19 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B20 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N12);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => HOLD0, A1 => UQVN_N6);
UQVB_B22 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B23 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => HOLD1, A1 => UQVN_N17);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => QI1);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => QI0);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => LD);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CS);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => DNUP);
UQVB_B29 : OR6
	PORT MAP (Z0 => UQVN_N17, A0 => LOAD1, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16);
UQVB_B30 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N13, A2 => UQVN_N12);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => LD);
UQVB_B32 : OR5
	PORT MAP (Z0 => UQVN_N24, A0 => LOAD2, A1 => UQVN_N26, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => CS);
UQVB_B34 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N30, A2 => UQVN_N31);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => DNUP);
UQVB_B36 : AND8
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N38, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => UQVN_N27, 
	A7 => UQVN_N31);
UQVB_B37 : AND8
	PORT MAP (Z0 => UQVN_N18, A0 => QI3, A1 => UQVN_N36, A2 => UQVN_N35, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N31);
UQVB_B38 : AND8
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N36, A2 => UQVN_N35, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N31);
UQVB_B39 : AND6
	PORT MAP (Z0 => UQVN_N20, A0 => QI3, A1 => QI2, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N31);
UQVB_B40 : AND8
	PORT MAP (Z0 => UQVN_N22, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => UQVN_N27, 
	A7 => UQVN_N31);
UQVB_B41 : AND7
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI0, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N27, A6 => UQVN_N31);
UQVB_B42 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N35, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N31);
UQVB_B43 : AND6
	PORT MAP (Z0 => UQVN_N29, A0 => QI3, A1 => QI2, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N31);
UQVB_B44 : AND6
	PORT MAP (Z0 => UQVN_N32, A0 => QI3, A1 => QI1, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N31);
UQVB_B45 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N31);
UQVB_B46 : OR6
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N21, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => UQVN_N28, A4 => UQVN_N29, A5 => UQVN_N32);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D3, A1 => LD, A2 => UQVN_N31);
UQVB_B48 : LXOR2
	PORT MAP (Z0 => UQVN_N25, A0 => HOLD3, A1 => UQVN_N33);
UQVB_B49 : LXOR2
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD2, A1 => UQVN_N24);
UQVB_B50 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => QI2);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => QI3);
UQVB_B53 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N25, CLK => CLK, CD => CD);
UQVB_B54 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N30, A2 => UQVN_N31);
END lattice_arch;
-- VHDL netlist for CDUD8
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDUD8 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END CDUD8;


ARCHITECTURE lattice_arch OF CDUD8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 HOLD0, HOLD1, HOLD2, HOLD3,
	 HOLD4, HOLD5, HOLD6, HOLD7,
	 LOAD0, LOAD1, LOAD2, LOAD4,
	 LOAD5, LOAD6, LOAD7, QI0,
	 QI1, QI2, QI3, QI4,
	 QI5, QI6, QI7, UQVN_N73,
	 UQVN_N74, UQVN_N75, UQVN_N76, UQVN_N77,
	 UQVN_N78, UQVN_N79, UQVN_N80 : std_logic;


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


BEGIN

UQVB_B1 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => QI0, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N4, A0 => LOAD0, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B3 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N11, A2 => UQVN_N10);
UQVB_B4 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => QI3, A1 => QI1, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B13 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N10);
UQVB_B14 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B15 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N10);
UQVB_B16 : LXOR2
	PORT MAP (Z0 => UQVN_N5, A0 => HOLD0, A1 => UQVN_N4);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N76, A1 => UQVN_N11, A2 => EN, 
	A3 => UQVN_N10);
UQVB_B18 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N75, A1 => UQVN_N74, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N10);
UQVB_B19 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => UQVN_N6, A0 => HOLD1, A1 => UQVN_N15);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N74, A0 => QI1);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N73, A0 => QI0);
UQVB_B23 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N76, A1 => QI0, A2 => UQVN_N11, 
	A3 => EN, A4 => UQVN_N12, A5 => UQVN_N10);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => LD);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B26 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => QI1, A1 => UQVN_N73, A2 => UQVN_N11, 
	A3 => EN, A4 => DNUP, A5 => UQVN_N10);
UQVB_B27 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N76, A1 => QI2, A2 => UQVN_N73, 
	A3 => UQVN_N11, A4 => EN, A5 => DNUP, A6 => UQVN_N10);
UQVB_B28 : AND7
	PORT MAP (Z0 => UQVN_N13, A0 => QI3, A1 => UQVN_N75, A2 => UQVN_N73, 
	A3 => UQVN_N11, A4 => EN, A5 => DNUP, A6 => UQVN_N10);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => DNUP);
UQVB_B30 : OR6
	PORT MAP (Z0 => UQVN_N15, A0 => LOAD1, A1 => UQVN_N7, A2 => UQVN_N8, 
	A3 => UQVN_N9, A4 => UQVN_N13, A5 => UQVN_N14);
UQVB_B31 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N11, A2 => UQVN_N10);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => LD);
UQVB_B33 : AND7
	PORT MAP (Z0 => UQVN_N17, A0 => QI2, A1 => UQVN_N74, A2 => UQVN_N73, 
	A3 => UQVN_N28, A4 => EN, A5 => DNUP, A6 => UQVN_N29);
UQVB_B34 : AND5
	PORT MAP (Z0 => UQVN_N18, A0 => QI3, A1 => QI2, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N29);
UQVB_B35 : OR5
	PORT MAP (Z0 => UQVN_N22, A0 => LOAD2, A1 => UQVN_N24, A2 => UQVN_N16, 
	A3 => UQVN_N17, A4 => UQVN_N18);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => CS);
UQVB_B37 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N28, A2 => UQVN_N29);
UQVB_B38 : AND5
	PORT MAP (Z0 => UQVN_N27, A0 => QI3, A1 => QI2, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N29);
UQVB_B39 : AND5
	PORT MAP (Z0 => UQVN_N30, A0 => QI3, A1 => QI1, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N29);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => DNUP);
UQVB_B41 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N29);
UQVB_B42 : AND7
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N76, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N28, A4 => EN, A5 => UQVN_N25, A6 => UQVN_N29);
UQVB_B43 : OR6
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N19, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N26, A4 => UQVN_N27, A5 => UQVN_N30);
UQVB_B44 : AND7
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => UQVN_N74, A2 => UQVN_N73, 
	A3 => UQVN_N28, A4 => EN, A5 => DNUP, A6 => UQVN_N29);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => D3, A1 => LD, A2 => UQVN_N29);
UQVB_B46 : AND7
	PORT MAP (Z0 => UQVN_N20, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N28, A4 => EN, A5 => UQVN_N25, A6 => UQVN_N29);
UQVB_B47 : AND6
	PORT MAP (Z0 => UQVN_N21, A0 => QI3, A1 => QI0, A2 => UQVN_N28, 
	A3 => EN, A4 => UQVN_N25, A5 => UQVN_N29);
UQVB_B48 : AND7
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N75, A1 => UQVN_N74, A2 => UQVN_N73, 
	A3 => UQVN_N28, A4 => EN, A5 => DNUP, A6 => UQVN_N29);
UQVB_B49 : LXOR2
	PORT MAP (Z0 => UQVN_N23, A0 => HOLD3, A1 => UQVN_N31);
UQVB_B50 : LXOR2
	PORT MAP (Z0 => UQVN_N32, A0 => HOLD2, A1 => UQVN_N22);
UQVB_B51 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N32, CLK => CLK, CD => CD);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N75, A0 => QI2);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N76, A0 => QI3);
UQVB_B54 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N23, CLK => CLK, CD => CD);
UQVB_B55 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N28, A2 => UQVN_N29);
UQVB_B56 : AND3
	PORT MAP (Z0 => LOAD4, A0 => D4, A1 => LD, A2 => UQVN_N40);
UQVB_B57 : AND9
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N80, A1 => QI3, A2 => UQVN_N75, 
	A3 => UQVN_N74, A4 => QI0, A5 => UQVN_N39, A6 => EN, 
	A7 => UQVN_N41, A8 => UQVN_N40);
UQVB_B58 : AND10
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N79, A1 => UQVN_N78, A2 => QI3, 
	A3 => UQVN_N75, A4 => UQVN_N74, A5 => QI0, A6 => UQVN_N39, 
	A7 => EN, A8 => UQVN_N41, A9 => UQVN_N40);
UQVB_B59 : AND9
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N80, A1 => UQVN_N76, A2 => UQVN_N75, 
	A3 => UQVN_N74, A4 => UQVN_N73, A5 => UQVN_N39, A6 => EN, 
	A7 => DNUP, A8 => UQVN_N40);
UQVB_B60 : AND10
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N79, A1 => UQVN_N78, A2 => UQVN_N76, 
	A3 => UQVN_N75, A4 => UQVN_N74, A5 => UQVN_N73, A6 => UQVN_N39, 
	A7 => EN, A8 => DNUP, A9 => UQVN_N40);
UQVB_B61 : OR7
	PORT MAP (Z0 => UQVN_N37, A0 => LOAD4, A1 => UQVN_N34, A2 => UQVN_N33, 
	A3 => UQVN_N35, A4 => UQVN_N36, A5 => UQVN_N42, A6 => UQVN_N43);
UQVB_B62 : LXOR2
	PORT MAP (Z0 => UQVN_N38, A0 => HOLD4, A1 => UQVN_N37);
UQVB_B63 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N38, CLK => CLK, CD => CD);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N77, A0 => QI4);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => LD);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CS);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => DNUP);
UQVB_B68 : AND3
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N39, A2 => UQVN_N40);
UQVB_B69 : AND6
	PORT MAP (Z0 => UQVN_N42, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N39, A4 => EN, A5 => UQVN_N40);
UQVB_B70 : AND6
	PORT MAP (Z0 => UQVN_N43, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N39, A4 => EN, A5 => UQVN_N40);
UQVB_B71 : AND3
	PORT MAP (Z0 => LOAD5, A0 => D5, A1 => LD, A2 => UQVN_N51);
UQVB_B72 : AND10
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N80, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N75, A4 => UQVN_N74, A5 => QI0, A6 => UQVN_N50, 
	A7 => EN, A8 => UQVN_N52, A9 => UQVN_N51);
UQVB_B73 : AND10
	PORT MAP (Z0 => UQVN_N44, A0 => QI5, A1 => UQVN_N77, A2 => UQVN_N76, 
	A3 => UQVN_N75, A4 => UQVN_N74, A5 => UQVN_N73, A6 => UQVN_N50, 
	A7 => EN, A8 => DNUP, A9 => UQVN_N51);
UQVB_B74 : AND11
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N80, A1 => QI6, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N75, A5 => UQVN_N74, A6 => UQVN_N73, 
	A7 => UQVN_N50, A8 => EN, A9 => DNUP, A10 => UQVN_N51);
UQVB_B75 : AND11
	PORT MAP (Z0 => UQVN_N49, A0 => QI7, A1 => UQVN_N79, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N75, A5 => UQVN_N74, A6 => UQVN_N73, 
	A7 => UQVN_N50, A8 => EN, A9 => DNUP, A10 => UQVN_N51);
UQVB_B76 : LXOR2
	PORT MAP (Z0 => UQVN_N46, A0 => HOLD5, A1 => UQVN_N45);
UQVB_B77 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N46, CLK => CLK, CD => CD);
UQVB_B78 : INV
	PORT MAP (ZN0 => UQVN_N78, A0 => QI5);
UQVB_B79 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => LD);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => CS);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => DNUP);
UQVB_B82 : AND3
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N50, A2 => UQVN_N51);
UQVB_B83 : AND5
	PORT MAP (Z0 => UQVN_N53, A0 => QI7, A1 => QI5, A2 => UQVN_N50, 
	A3 => EN, A4 => UQVN_N51);
UQVB_B84 : OR6
	PORT MAP (Z0 => UQVN_N45, A0 => LOAD5, A1 => UQVN_N47, A2 => UQVN_N44, 
	A3 => UQVN_N48, A4 => UQVN_N49, A5 => UQVN_N53);
UQVB_B85 : AND3
	PORT MAP (Z0 => LOAD6, A0 => D6, A1 => LD, A2 => UQVN_N60);
UQVB_B86 : AND11
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N80, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N75, A5 => UQVN_N74, A6 => QI0, 
	A7 => UQVN_N59, A8 => EN, A9 => UQVN_N61, A10 => UQVN_N60);
UQVB_B87 : AND11
	PORT MAP (Z0 => UQVN_N54, A0 => QI7, A1 => UQVN_N78, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N75, A5 => UQVN_N74, A6 => UQVN_N73, 
	A7 => UQVN_N59, A8 => EN, A9 => DNUP, A10 => UQVN_N60);
UQVB_B88 : AND11
	PORT MAP (Z0 => UQVN_N58, A0 => QI6, A1 => UQVN_N78, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N75, A5 => UQVN_N74, A6 => UQVN_N73, 
	A7 => UQVN_N59, A8 => EN, A9 => DNUP, A10 => UQVN_N60);
UQVB_B89 : LXOR2
	PORT MAP (Z0 => UQVN_N56, A0 => HOLD6, A1 => UQVN_N55);
UQVB_B90 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N56, CLK => CLK, CD => CD);
UQVB_B91 : INV
	PORT MAP (ZN0 => UQVN_N79, A0 => QI6);
UQVB_B92 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => LD);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N60, A0 => CS);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N61, A0 => DNUP);
UQVB_B95 : AND3
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N59, A2 => UQVN_N60);
UQVB_B96 : AND5
	PORT MAP (Z0 => UQVN_N62, A0 => QI7, A1 => QI6, A2 => UQVN_N59, 
	A3 => EN, A4 => UQVN_N60);
UQVB_B97 : OR5
	PORT MAP (Z0 => UQVN_N55, A0 => LOAD6, A1 => UQVN_N57, A2 => UQVN_N54, 
	A3 => UQVN_N58, A4 => UQVN_N62);
UQVB_B98 : AND3
	PORT MAP (Z0 => LOAD7, A0 => D7, A1 => LD, A2 => UQVN_N70);
UQVB_B99 : AND11
	PORT MAP (Z0 => UQVN_N64, A0 => QI6, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N75, A5 => UQVN_N74, A6 => QI0, 
	A7 => UQVN_N69, A8 => EN, A9 => UQVN_N71, A10 => UQVN_N70);
UQVB_B100 : AND10
	PORT MAP (Z0 => UQVN_N63, A0 => QI7, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N75, A4 => UQVN_N74, A5 => QI0, A6 => UQVN_N69, 
	A7 => EN, A8 => UQVN_N71, A9 => UQVN_N70);
UQVB_B101 : AND11
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N79, A1 => UQVN_N78, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N75, A5 => UQVN_N74, A6 => UQVN_N73, 
	A7 => UQVN_N69, A8 => EN, A9 => DNUP, A10 => UQVN_N70);
UQVB_B102 : LXOR2
	PORT MAP (Z0 => UQVN_N68, A0 => HOLD7, A1 => UQVN_N67);
UQVB_B103 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N68, CLK => CLK, CD => CD);
UQVB_B104 : INV
	PORT MAP (ZN0 => UQVN_N80, A0 => QI7);
UQVB_B105 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => LD);
UQVB_B106 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => DNUP);
UQVB_B107 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => CS);
UQVB_B108 : AND3
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N69, A2 => UQVN_N70);
UQVB_B109 : AND5
	PORT MAP (Z0 => UQVN_N66, A0 => QI7, A1 => QI6, A2 => UQVN_N69, 
	A3 => EN, A4 => UQVN_N70);
UQVB_B110 : AND5
	PORT MAP (Z0 => UQVN_N72, A0 => QI7, A1 => QI5, A2 => UQVN_N69, 
	A3 => EN, A4 => UQVN_N70);
UQVB_B111 : OR6
	PORT MAP (Z0 => UQVN_N67, A0 => LOAD7, A1 => UQVN_N64, A2 => UQVN_N63, 
	A3 => UQVN_N65, A4 => UQVN_N66, A5 => UQVN_N72);
END lattice_arch;
-- VHDL netlist for CDUD8C
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CDUD8C IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic;
        CAO : OUT std_logic
    );
END CDUD8C;


ARCHITECTURE lattice_arch OF CDUD8C IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, HOLD0, HOLD1,
	 HOLD2, HOLD3, HOLD4, HOLD5,
	 HOLD6, HOLD7, LOAD0, LOAD1,
	 LOAD2, LOAD4, LOAD5, LOAD6,
	 LOAD7, QI0, QI1, QI2,
	 QI3, QI4, QI5, QI6,
	 QI7, UQVN_N75, UQVN_N76, UQVN_N77,
	 UQVN_N78, UQVN_N79, UQVN_N80, UQVN_N81,
	 UQVN_N82 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT AND10
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND10 use  entity  lat_vhd.AND10(lattice_arch);


  COMPONENT AND12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND12 use  entity  lat_vhd.AND12(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N6, A0 => LOAD0, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B2 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N13, A2 => UQVN_N12);
UQVB_B3 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N78, A1 => UQVN_N13, A2 => EN, 
	A3 => CAI, A4 => UQVN_N12);
UQVB_B4 : AND6
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N77, A1 => UQVN_N76, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N12);
UQVB_B5 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => QI3, A1 => QI0, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N12);
UQVB_B6 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N78, A1 => QI0, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N14, A6 => UQVN_N12);
UQVB_B7 : AND7
	PORT MAP (Z0 => UQVN_N10, A0 => QI1, A1 => UQVN_N75, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => DNUP, A6 => UQVN_N12);
UQVB_B8 : AND8
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N78, A1 => QI2, A2 => UQVN_N75, 
	A3 => UQVN_N13, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N12);
UQVB_B9 : AND8
	PORT MAP (Z0 => UQVN_N15, A0 => QI3, A1 => UQVN_N77, A2 => UQVN_N75, 
	A3 => UQVN_N13, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N12);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI1, A2 => UQVN_N13, 
	A3 => EN, A4 => CAI, A5 => UQVN_N12);
UQVB_B11 : AND11
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N82, A1 => UQVN_N81, A2 => UQVN_N80, 
	A3 => UQVN_N79, A4 => UQVN_N78, A5 => UQVN_N77, A6 => UQVN_N76, 
	A7 => UQVN_N75, A8 => EN, A9 => CAI, A10 => DNUP);
UQVB_B12 : AND11
	PORT MAP (Z0 => UQVN_N4, A0 => QI7, A1 => UQVN_N81, A2 => UQVN_N80, 
	A3 => QI4, A4 => QI3, A5 => UQVN_N77, A6 => UQVN_N76, 
	A7 => QI0, A8 => EN, A9 => CAI, A10 => UQVN_N14);
UQVB_B13 : OR2
	PORT MAP (Z0 => CAO, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q4, A0 => QI4);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q5, A0 => QI5);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q6, A0 => QI6);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q7, A0 => QI7);
UQVB_B22 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N12);
UQVB_B23 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B24 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N12);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => UQVN_N7, A0 => HOLD0, A1 => UQVN_N6);
UQVB_B26 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B27 : LXOR2
	PORT MAP (Z0 => UQVN_N8, A0 => HOLD1, A1 => UQVN_N17);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N76, A0 => QI1);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N75, A0 => QI0);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => LD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CS);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => DNUP);
UQVB_B33 : OR6
	PORT MAP (Z0 => UQVN_N17, A0 => LOAD1, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16);
UQVB_B34 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N13, A2 => UQVN_N12);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => LD);
UQVB_B36 : OR5
	PORT MAP (Z0 => UQVN_N24, A0 => LOAD2, A1 => UQVN_N26, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => CS);
UQVB_B38 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N30, A2 => UQVN_N31);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => DNUP);
UQVB_B40 : AND8
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N78, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => UQVN_N27, 
	A7 => UQVN_N31);
UQVB_B41 : AND8
	PORT MAP (Z0 => UQVN_N18, A0 => QI3, A1 => UQVN_N76, A2 => UQVN_N75, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N31);
UQVB_B42 : AND8
	PORT MAP (Z0 => UQVN_N19, A0 => QI2, A1 => UQVN_N76, A2 => UQVN_N75, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N31);
UQVB_B43 : AND6
	PORT MAP (Z0 => UQVN_N20, A0 => QI3, A1 => QI2, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N31);
UQVB_B44 : AND8
	PORT MAP (Z0 => UQVN_N22, A0 => QI2, A1 => QI1, A2 => QI0, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => UQVN_N27, 
	A7 => UQVN_N31);
UQVB_B45 : AND7
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI0, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N27, A6 => UQVN_N31);
UQVB_B46 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N77, A1 => UQVN_N76, A2 => UQVN_N75, 
	A3 => UQVN_N30, A4 => EN, A5 => CAI, A6 => DNUP, 
	A7 => UQVN_N31);
UQVB_B47 : AND6
	PORT MAP (Z0 => UQVN_N29, A0 => QI3, A1 => QI2, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N31);
UQVB_B48 : AND6
	PORT MAP (Z0 => UQVN_N32, A0 => QI3, A1 => QI1, A2 => UQVN_N30, 
	A3 => EN, A4 => CAI, A5 => UQVN_N31);
UQVB_B49 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N31);
UQVB_B50 : OR6
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N21, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => UQVN_N28, A4 => UQVN_N29, A5 => UQVN_N32);
UQVB_B51 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D3, A1 => LD, A2 => UQVN_N31);
UQVB_B52 : LXOR2
	PORT MAP (Z0 => UQVN_N25, A0 => HOLD3, A1 => UQVN_N33);
UQVB_B53 : LXOR2
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD2, A1 => UQVN_N24);
UQVB_B54 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N77, A0 => QI2);
UQVB_B56 : INV
	PORT MAP (ZN0 => UQVN_N78, A0 => QI3);
UQVB_B57 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N25, CLK => CLK, CD => CD);
UQVB_B58 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N30, A2 => UQVN_N31);
UQVB_B59 : AND3
	PORT MAP (Z0 => LOAD4, A0 => D4, A1 => LD, A2 => UQVN_N42);
UQVB_B60 : OR7
	PORT MAP (Z0 => UQVN_N39, A0 => LOAD4, A1 => UQVN_N36, A2 => UQVN_N35, 
	A3 => UQVN_N37, A4 => UQVN_N38, A5 => UQVN_N44, A6 => UQVN_N45);
UQVB_B61 : LXOR2
	PORT MAP (Z0 => UQVN_N40, A0 => HOLD4, A1 => UQVN_N39);
UQVB_B62 : FD21
	PORT MAP (Q0 => QI4, D0 => UQVN_N40, CLK => CLK, CD => CD);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N79, A0 => QI4);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => LD);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => CS);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => DNUP);
UQVB_B67 : AND3
	PORT MAP (Z0 => HOLD4, A0 => QI4, A1 => UQVN_N41, A2 => UQVN_N42);
UQVB_B68 : AND10
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N82, A1 => QI3, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => QI0, A5 => UQVN_N41, A6 => EN, 
	A7 => CAI, A8 => UQVN_N43, A9 => UQVN_N42);
UQVB_B69 : AND11
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N81, A1 => UQVN_N80, A2 => QI3, 
	A3 => UQVN_N77, A4 => UQVN_N76, A5 => QI0, A6 => UQVN_N41, 
	A7 => EN, A8 => CAI, A9 => UQVN_N43, A10 => UQVN_N42);
UQVB_B70 : AND10
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N82, A1 => UQVN_N78, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N75, A5 => UQVN_N41, A6 => EN, 
	A7 => CAI, A8 => DNUP, A9 => UQVN_N42);
UQVB_B71 : AND11
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N81, A1 => UQVN_N80, A2 => UQVN_N78, 
	A3 => UQVN_N77, A4 => UQVN_N76, A5 => UQVN_N75, A6 => UQVN_N41, 
	A7 => EN, A8 => CAI, A9 => DNUP, A10 => UQVN_N42);
UQVB_B72 : AND7
	PORT MAP (Z0 => UQVN_N44, A0 => QI7, A1 => QI6, A2 => QI4, 
	A3 => UQVN_N41, A4 => EN, A5 => CAI, A6 => UQVN_N42);
UQVB_B73 : AND7
	PORT MAP (Z0 => UQVN_N45, A0 => QI7, A1 => QI5, A2 => QI4, 
	A3 => UQVN_N41, A4 => EN, A5 => CAI, A6 => UQVN_N42);
UQVB_B74 : AND3
	PORT MAP (Z0 => LOAD5, A0 => D5, A1 => LD, A2 => UQVN_N53);
UQVB_B75 : LXOR2
	PORT MAP (Z0 => UQVN_N48, A0 => HOLD5, A1 => UQVN_N47);
UQVB_B76 : FD21
	PORT MAP (Q0 => QI5, D0 => UQVN_N48, CLK => CLK, CD => CD);
UQVB_B77 : INV
	PORT MAP (ZN0 => UQVN_N80, A0 => QI5);
UQVB_B78 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => LD);
UQVB_B79 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => CS);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => DNUP);
UQVB_B81 : AND3
	PORT MAP (Z0 => HOLD5, A0 => QI5, A1 => UQVN_N52, A2 => UQVN_N53);
UQVB_B82 : OR6
	PORT MAP (Z0 => UQVN_N47, A0 => LOAD5, A1 => UQVN_N49, A2 => UQVN_N46, 
	A3 => UQVN_N50, A4 => UQVN_N51, A5 => UQVN_N55);
UQVB_B83 : AND11
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N82, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N77, A4 => UQVN_N76, A5 => QI0, A6 => UQVN_N52, 
	A7 => EN, A8 => CAI, A9 => UQVN_N54, A10 => UQVN_N53);
UQVB_B84 : AND11
	PORT MAP (Z0 => UQVN_N46, A0 => QI5, A1 => UQVN_N79, A2 => UQVN_N78, 
	A3 => UQVN_N77, A4 => UQVN_N76, A5 => UQVN_N75, A6 => UQVN_N52, 
	A7 => EN, A8 => CAI, A9 => DNUP, A10 => UQVN_N53);
UQVB_B85 : AND12
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N82, A1 => QI6, A2 => UQVN_N79, 
	A3 => UQVN_N78, A4 => UQVN_N77, A5 => UQVN_N76, A6 => UQVN_N75, 
	A7 => UQVN_N52, A8 => EN, A9 => CAI, A10 => DNUP, 
	A11 => UQVN_N53);
UQVB_B86 : AND12
	PORT MAP (Z0 => UQVN_N51, A0 => QI7, A1 => UQVN_N81, A2 => UQVN_N79, 
	A3 => UQVN_N78, A4 => UQVN_N77, A5 => UQVN_N76, A6 => UQVN_N75, 
	A7 => UQVN_N52, A8 => EN, A9 => CAI, A10 => DNUP, 
	A11 => UQVN_N53);
UQVB_B87 : AND6
	PORT MAP (Z0 => UQVN_N55, A0 => QI7, A1 => QI5, A2 => UQVN_N52, 
	A3 => EN, A4 => CAI, A5 => UQVN_N53);
UQVB_B88 : AND3
	PORT MAP (Z0 => LOAD6, A0 => D6, A1 => LD, A2 => UQVN_N62);
UQVB_B89 : LXOR2
	PORT MAP (Z0 => UQVN_N58, A0 => HOLD6, A1 => UQVN_N57);
UQVB_B90 : FD21
	PORT MAP (Q0 => QI6, D0 => UQVN_N58, CLK => CLK, CD => CD);
UQVB_B91 : INV
	PORT MAP (ZN0 => UQVN_N81, A0 => QI6);
UQVB_B92 : INV
	PORT MAP (ZN0 => UQVN_N61, A0 => LD);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => CS);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N63, A0 => DNUP);
UQVB_B95 : AND3
	PORT MAP (Z0 => HOLD6, A0 => QI6, A1 => UQVN_N61, A2 => UQVN_N62);
UQVB_B96 : OR5
	PORT MAP (Z0 => UQVN_N57, A0 => LOAD6, A1 => UQVN_N59, A2 => UQVN_N56, 
	A3 => UQVN_N60, A4 => UQVN_N64);
UQVB_B97 : AND12
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N82, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N77, A5 => UQVN_N76, A6 => QI0, 
	A7 => UQVN_N61, A8 => EN, A9 => CAI, A10 => UQVN_N63, 
	A11 => UQVN_N62);
UQVB_B98 : AND12
	PORT MAP (Z0 => UQVN_N56, A0 => QI7, A1 => UQVN_N80, A2 => UQVN_N79, 
	A3 => UQVN_N78, A4 => UQVN_N77, A5 => UQVN_N76, A6 => UQVN_N75, 
	A7 => UQVN_N61, A8 => EN, A9 => CAI, A10 => DNUP, 
	A11 => UQVN_N62);
UQVB_B99 : AND12
	PORT MAP (Z0 => UQVN_N60, A0 => QI6, A1 => UQVN_N80, A2 => UQVN_N79, 
	A3 => UQVN_N78, A4 => UQVN_N77, A5 => UQVN_N76, A6 => UQVN_N75, 
	A7 => UQVN_N61, A8 => EN, A9 => CAI, A10 => DNUP, 
	A11 => UQVN_N62);
UQVB_B100 : AND6
	PORT MAP (Z0 => UQVN_N64, A0 => QI7, A1 => QI6, A2 => UQVN_N61, 
	A3 => EN, A4 => CAI, A5 => UQVN_N62);
UQVB_B101 : AND3
	PORT MAP (Z0 => LOAD7, A0 => D7, A1 => LD, A2 => UQVN_N72);
UQVB_B102 : LXOR2
	PORT MAP (Z0 => UQVN_N70, A0 => HOLD7, A1 => UQVN_N69);
UQVB_B103 : FD21
	PORT MAP (Q0 => QI7, D0 => UQVN_N70, CLK => CLK, CD => CD);
UQVB_B104 : INV
	PORT MAP (ZN0 => UQVN_N82, A0 => QI7);
UQVB_B105 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => LD);
UQVB_B106 : INV
	PORT MAP (ZN0 => UQVN_N73, A0 => DNUP);
UQVB_B107 : INV
	PORT MAP (ZN0 => UQVN_N72, A0 => CS);
UQVB_B108 : AND3
	PORT MAP (Z0 => HOLD7, A0 => QI7, A1 => UQVN_N71, A2 => UQVN_N72);
UQVB_B109 : OR6
	PORT MAP (Z0 => UQVN_N69, A0 => LOAD7, A1 => UQVN_N66, A2 => UQVN_N65, 
	A3 => UQVN_N67, A4 => UQVN_N68, A5 => UQVN_N74);
UQVB_B110 : AND12
	PORT MAP (Z0 => UQVN_N66, A0 => QI6, A1 => QI5, A2 => QI4, 
	A3 => QI3, A4 => UQVN_N77, A5 => UQVN_N76, A6 => QI0, 
	A7 => UQVN_N71, A8 => EN, A9 => CAI, A10 => UQVN_N73, 
	A11 => UQVN_N72);
UQVB_B111 : AND11
	PORT MAP (Z0 => UQVN_N65, A0 => QI7, A1 => QI4, A2 => QI3, 
	A3 => UQVN_N77, A4 => UQVN_N76, A5 => QI0, A6 => UQVN_N71, 
	A7 => EN, A8 => CAI, A9 => UQVN_N73, A10 => UQVN_N72);
UQVB_B112 : AND12
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N81, A1 => UQVN_N80, A2 => UQVN_N79, 
	A3 => UQVN_N78, A4 => UQVN_N77, A5 => UQVN_N76, A6 => UQVN_N75, 
	A7 => UQVN_N71, A8 => EN, A9 => CAI, A10 => DNUP, 
	A11 => UQVN_N72);
UQVB_B113 : AND6
	PORT MAP (Z0 => UQVN_N68, A0 => QI7, A1 => QI6, A2 => UQVN_N71, 
	A3 => EN, A4 => CAI, A5 => UQVN_N72);
UQVB_B114 : AND6
	PORT MAP (Z0 => UQVN_N74, A0 => QI7, A1 => QI5, A2 => UQVN_N71, 
	A3 => EN, A4 => CAI, A5 => UQVN_N72);
END lattice_arch;
-- VHDL netlist for CGD14
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CGD14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CGD14;


ARCHITECTURE lattice_arch OF CGD14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, HOLD0, HOLD1, HOLD2,
	 HOLD3, LOAD0, LOAD1, LOAD2,
	 LOAD3, QI0, QI1, QI2,
	 QI3, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25 : std_logic;


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => UQVN_N24, A2 => QI0, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B2 : OR7
	PORT MAP (Z0 => UQVN_N9, A0 => HOLD0, A1 => LOAD0, A2 => UQVN_N1, 
	A3 => UQVN_N10, A4 => UQVN_N2, A5 => UQVN_N4, A6 => PS);
UQVB_B3 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N8, A2 => UQVN_N3);
UQVB_B4 : AND2
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD);
UQVB_B5 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N25, A1 => UQVN_N24, A2 => QI1, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N25, A1 => QI2, A2 => UQVN_N23, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI2, A2 => QI1, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B9 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N8, A2 => UQVN_N3);
UQVB_B10 : AND2
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N25, A1 => QI2, A2 => QI0, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B12 : OR6
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD1, A1 => LOAD1, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N7, A5 => PS);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => LD);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => EN);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B19 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B20 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI1);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => QI0);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => QI1, A1 => UQVN_N22, A2 => UQVN_N8, 
	A3 => EN);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => LD);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => EN);
UQVB_B26 : OR6
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD3, A1 => LOAD3, A2 => UQVN_N12, 
	A3 => UQVN_N20, A4 => UQVN_N21, A5 => PS);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI3);
UQVB_B28 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI3, A1 => QI1, A2 => UQVN_N22, 
	A3 => UQVN_N19, A4 => EN);
UQVB_B29 : AND2
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI2);
UQVB_B31 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => QI2, A1 => UQVN_N23, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B32 : OR6
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD2, A1 => LOAD2, A2 => UQVN_N16, 
	A3 => UQVN_N15, A4 => UQVN_N14, A5 => PS);
UQVB_B33 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B34 : AND2
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N22, 
	A3 => UQVN_N19, A4 => EN);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => QI2, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B39 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B40 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N17, CLK => CLK, CD => CD);
UQVB_B41 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N13, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CGD24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CGD24 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CGD24;


ARCHITECTURE lattice_arch OF CGD24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, HOLD0,
	 HOLD1, HOLD2, HOLD3, LOAD0,
	 LOAD1, LOAD2, LOAD3, QI0,
	 QI1, QI2, QI3, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


BEGIN

UQVB_B1 : OR7
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD0, A1 => LOAD0, A2 => UQVN_N1, 
	A3 => UQVN_N11, A4 => UQVN_N7, A5 => UQVN_N8, A6 => PS);
UQVB_B2 : OR6
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD1, A1 => LOAD1, A2 => UQVN_N4, 
	A3 => UQVN_N3, A4 => UQVN_N5, A5 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => LD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N6, A2 => UQVN_N2, 
	A3 => UQVN_N9);
UQVB_B6 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N9);
UQVB_B7 : AND6
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N27, A1 => UQVN_N26, A2 => QI1, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B8 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N27, A1 => QI2, A2 => UQVN_N25, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI2, A2 => QI1, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => UQVN_N26, A2 => UQVN_N25, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B11 : AND4
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N6, A2 => UQVN_N2, 
	A3 => UQVN_N9);
UQVB_B12 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N9);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI1, A1 => UQVN_N24, A2 => UQVN_N6, 
	A3 => EN, A4 => UQVN_N9);
UQVB_B14 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N27, A1 => QI2, A2 => QI0, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => UQVN_N26, A2 => QI0, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => CS);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B21 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N10, CLK => CLK);
UQVB_B22 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N12, CLK => CLK);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI0);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => LD);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => EN);
UQVB_B27 : AND4
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N14);
UQVB_B28 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N14);
UQVB_B29 : AND6
	PORT MAP (Z0 => UQVN_N18, A0 => QI3, A1 => QI1, A2 => UQVN_N24, 
	A3 => UQVN_N21, A4 => EN, A5 => UQVN_N14);
UQVB_B30 : AND5
	PORT MAP (Z0 => UQVN_N17, A0 => QI2, A1 => UQVN_N25, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B31 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI2, A1 => QI0, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B32 : AND4
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N14);
UQVB_B33 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N14);
UQVB_B34 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N21, A4 => EN, A5 => UQVN_N14);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => QI0, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B36 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI1, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => CS);
UQVB_B38 : OR6
	PORT MAP (Z0 => UQVN_N15, A0 => HOLD3, A1 => LOAD3, A2 => UQVN_N13, 
	A3 => UQVN_N22, A4 => UQVN_N23, A5 => PS);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B41 : OR6
	PORT MAP (Z0 => UQVN_N19, A0 => HOLD2, A1 => LOAD2, A2 => UQVN_N18, 
	A3 => UQVN_N17, A4 => UQVN_N16, A5 => PS);
UQVB_B42 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N19, CLK => CLK);
UQVB_B43 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N15, CLK => CLK);
END lattice_arch;
-- VHDL netlist for CGU14
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CGU14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CGU14;


ARCHITECTURE lattice_arch OF CGU14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, HOLD0, HOLD1, HOLD2,
	 HOLD3, LOAD0, LOAD1, LOAD2,
	 LOAD3, QI0, QI1, QI2,
	 QI3, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25 : std_logic;


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI2, A2 => QI0, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B2 : OR7
	PORT MAP (Z0 => UQVN_N9, A0 => HOLD0, A1 => LOAD0, A2 => UQVN_N1, 
	A3 => UQVN_N10, A4 => UQVN_N2, A5 => UQVN_N4, A6 => PS);
UQVB_B3 : AND3
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N8, A2 => UQVN_N3);
UQVB_B4 : AND2
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD);
UQVB_B5 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N25, A1 => QI2, A2 => QI1, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => QI3, A1 => QI2, A2 => UQVN_N23, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => UQVN_N24, A2 => QI1, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B9 : AND3
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N8, A2 => UQVN_N3);
UQVB_B10 : AND2
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N25, A1 => UQVN_N24, A2 => QI0, 
	A3 => UQVN_N8, A4 => EN);
UQVB_B12 : OR6
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD1, A1 => LOAD1, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N7, A5 => PS);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => LD);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => EN);
UQVB_B15 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B19 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N9, CLK => CLK, CD => CD);
UQVB_B20 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => QI1);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => QI0);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => QI1, A1 => UQVN_N22, A2 => UQVN_N8, 
	A3 => EN);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => LD);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => EN);
UQVB_B26 : OR6
	PORT MAP (Z0 => UQVN_N13, A0 => HOLD3, A1 => LOAD3, A2 => UQVN_N12, 
	A3 => UQVN_N20, A4 => UQVN_N21, A5 => PS);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI3);
UQVB_B28 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N25, A1 => QI1, A2 => UQVN_N22, 
	A3 => UQVN_N19, A4 => EN);
UQVB_B29 : AND2
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI2);
UQVB_B31 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => QI2, A1 => UQVN_N23, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B32 : OR6
	PORT MAP (Z0 => UQVN_N17, A0 => HOLD2, A1 => LOAD2, A2 => UQVN_N16, 
	A3 => UQVN_N15, A4 => UQVN_N14, A5 => PS);
UQVB_B33 : AND3
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B34 : AND2
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => QI2, A1 => UQVN_N23, A2 => UQVN_N22, 
	A3 => UQVN_N19, A4 => EN);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => QI3, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => QI3, A1 => QI1, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => QI2, A1 => QI0, A2 => UQVN_N19, 
	A3 => EN);
UQVB_B39 : AND3
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B40 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N17, CLK => CLK, CD => CD);
UQVB_B41 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N13, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CGU24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CGU24 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CGU24;


ARCHITECTURE lattice_arch OF CGU24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, HOLD0,
	 HOLD1, HOLD2, HOLD3, LOAD0,
	 LOAD1, LOAD2, LOAD3, QI0,
	 QI1, QI2, QI3, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27 : std_logic;


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


BEGIN

UQVB_B1 : OR7
	PORT MAP (Z0 => UQVN_N10, A0 => HOLD0, A1 => LOAD0, A2 => UQVN_N1, 
	A3 => UQVN_N11, A4 => UQVN_N7, A5 => UQVN_N8, A6 => PS);
UQVB_B2 : OR6
	PORT MAP (Z0 => UQVN_N12, A0 => HOLD1, A1 => LOAD1, A2 => UQVN_N4, 
	A3 => UQVN_N3, A4 => UQVN_N5, A5 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => LD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N6, A2 => UQVN_N2, 
	A3 => UQVN_N9);
UQVB_B6 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N9);
UQVB_B7 : AND6
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N25, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B8 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N27, A1 => QI2, A2 => QI1, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI2, A2 => UQVN_N25, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => QI3, A1 => UQVN_N26, A2 => QI1, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B11 : AND4
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N6, A2 => UQVN_N2, 
	A3 => UQVN_N9);
UQVB_B12 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N9);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => QI1, A1 => UQVN_N24, A2 => UQVN_N6, 
	A3 => EN, A4 => UQVN_N9);
UQVB_B14 : AND6
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N27, A1 => UQVN_N26, A2 => QI0, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => QI2, A2 => QI0, 
	A3 => UQVN_N6, A4 => EN, A5 => UQVN_N9);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => CS);
UQVB_B17 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B21 : FD11
	PORT MAP (Q0 => QI0, D0 => UQVN_N10, CLK => CLK);
UQVB_B22 : FD11
	PORT MAP (Q0 => QI1, D0 => UQVN_N12, CLK => CLK);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => QI1);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => QI0);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => LD);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => EN);
UQVB_B27 : AND4
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N14);
UQVB_B28 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N14);
UQVB_B29 : AND6
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N27, A1 => QI1, A2 => UQVN_N24, 
	A3 => UQVN_N21, A4 => EN, A5 => UQVN_N14);
UQVB_B30 : AND5
	PORT MAP (Z0 => UQVN_N17, A0 => QI2, A1 => UQVN_N25, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B31 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => QI2, A1 => QI0, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B32 : AND4
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N21, A2 => UQVN_N20, 
	A3 => UQVN_N14);
UQVB_B33 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N14);
UQVB_B34 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => QI2, A1 => UQVN_N25, A2 => UQVN_N24, 
	A3 => UQVN_N21, A4 => EN, A5 => UQVN_N14);
UQVB_B35 : AND5
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => QI0, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B36 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => QI3, A1 => QI1, A2 => UQVN_N21, 
	A3 => EN, A4 => UQVN_N14);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => CS);
UQVB_B38 : OR6
	PORT MAP (Z0 => UQVN_N15, A0 => HOLD3, A1 => LOAD3, A2 => UQVN_N13, 
	A3 => UQVN_N22, A4 => UQVN_N23, A5 => PS);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => QI3);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => QI2);
UQVB_B41 : OR6
	PORT MAP (Z0 => UQVN_N19, A0 => HOLD2, A1 => LOAD2, A2 => UQVN_N18, 
	A3 => UQVN_N17, A4 => UQVN_N16, A5 => PS);
UQVB_B42 : FD11
	PORT MAP (Q0 => QI2, D0 => UQVN_N19, CLK => CLK);
UQVB_B43 : FD11
	PORT MAP (Q0 => QI3, D0 => UQVN_N15, CLK => CLK);
END lattice_arch;
-- VHDL netlist for CGUD4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CGUD4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        DNUP : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END CGUD4;


ARCHITECTURE lattice_arch OF CGUD4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, HOLD0, HOLD1, HOLD2,
	 HOLD3, LOAD0, LOAD1, LOAD2,
	 LOAD3, QI0, QI1, QI2,
	 QI3, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45 : std_logic;


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : OR7
	PORT MAP (Z0 => UQVN_N11, A0 => HOLD0, A1 => LOAD0, A2 => UQVN_N1, 
	A3 => UQVN_N15, A4 => UQVN_N4, A5 => UQVN_N5, A6 => PS);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => EN);
UQVB_B3 : AND4
	PORT MAP (Z0 => HOLD0, A0 => QI0, A1 => UQVN_N3, A2 => UQVN_N2, 
	A3 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => LOAD0, A0 => D0, A1 => LD, A2 => UQVN_N6);
UQVB_B5 : AND7
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N45, A1 => UQVN_N44, A2 => UQVN_N43, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => UQVN_N14);
UQVB_B6 : AND7
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N45, A1 => QI2, A2 => QI1, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => UQVN_N14);
UQVB_B7 : AND7
	PORT MAP (Z0 => UQVN_N4, A0 => QI3, A1 => QI2, A2 => UQVN_N43, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => UQVN_N14);
UQVB_B8 : AND7
	PORT MAP (Z0 => UQVN_N5, A0 => QI3, A1 => UQVN_N44, A2 => QI1, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => UQVN_N14);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => LD);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => CS);
UQVB_B11 : AND7
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N45, A1 => UQVN_N44, A2 => QI1, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => DNUP);
UQVB_B12 : AND7
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N45, A1 => QI2, A2 => UQVN_N43, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => DNUP);
UQVB_B13 : AND7
	PORT MAP (Z0 => UQVN_N7, A0 => QI3, A1 => QI2, A2 => QI1, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => DNUP);
UQVB_B14 : AND7
	PORT MAP (Z0 => UQVN_N9, A0 => QI3, A1 => UQVN_N44, A2 => UQVN_N43, 
	A3 => UQVN_N3, A4 => EN, A5 => UQVN_N6, A6 => DNUP);
UQVB_B15 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N10, A1 => UQVN_N8, A2 => UQVN_N7, 
	A3 => UQVN_N9);
UQVB_B16 : OR2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => DNUP);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q3, A0 => QI3);
UQVB_B19 : BUF
	PORT MAP (Z0 => Q2, A0 => QI2);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q1, A0 => QI1);
UQVB_B21 : BUF
	PORT MAP (Z0 => Q0, A0 => QI0);
UQVB_B22 : FD21
	PORT MAP (Q0 => QI0, D0 => UQVN_N13, CLK => CLK, CD => CD);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => QI0);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => DNUP);
UQVB_B25 : FD21
	PORT MAP (Q0 => QI1, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => QI1);
UQVB_B27 : AND5
	PORT MAP (Z0 => UQVN_N18, A0 => QI1, A1 => UQVN_N42, A2 => UQVN_N16, 
	A3 => EN, A4 => UQVN_N19);
UQVB_B28 : AND4
	PORT MAP (Z0 => HOLD1, A0 => QI1, A1 => UQVN_N16, A2 => UQVN_N23, 
	A3 => UQVN_N19);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => EN);
UQVB_B30 : AND3
	PORT MAP (Z0 => LOAD1, A0 => D1, A1 => LD, A2 => UQVN_N19);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => CS);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => LD);
UQVB_B33 : AND7
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N45, A1 => UQVN_N44, A2 => QI0, 
	A3 => UQVN_N16, A4 => EN, A5 => UQVN_N19, A6 => UQVN_N27);
UQVB_B34 : AND7
	PORT MAP (Z0 => UQVN_N20, A0 => QI3, A1 => QI2, A2 => QI0, 
	A3 => UQVN_N16, A4 => EN, A5 => UQVN_N19, A6 => UQVN_N27);
UQVB_B35 : OR4
	PORT MAP (Z0 => UQVN_N24, A0 => HOLD1, A1 => LOAD1, A2 => PS, 
	A3 => UQVN_N18);
UQVB_B36 : AND7
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N45, A1 => QI2, A2 => QI0, 
	A3 => UQVN_N16, A4 => EN, A5 => UQVN_N19, A6 => DNUP);
UQVB_B37 : AND7
	PORT MAP (Z0 => UQVN_N22, A0 => QI3, A1 => UQVN_N44, A2 => QI0, 
	A3 => UQVN_N16, A4 => EN, A5 => UQVN_N19, A6 => DNUP);
UQVB_B38 : OR4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N17, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N22);
UQVB_B39 : OR2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N24, A1 => UQVN_N25);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => EN);
UQVB_B41 : AND4
	PORT MAP (Z0 => HOLD2, A0 => QI2, A1 => UQVN_N41, A2 => UQVN_N40, 
	A3 => UQVN_N28);
UQVB_B42 : AND3
	PORT MAP (Z0 => LOAD2, A0 => D2, A1 => LD, A2 => UQVN_N28);
UQVB_B43 : AND5
	PORT MAP (Z0 => UQVN_N37, A0 => QI2, A1 => UQVN_N43, A2 => UQVN_N41, 
	A3 => EN, A4 => UQVN_N28);
UQVB_B44 : AND5
	PORT MAP (Z0 => UQVN_N36, A0 => QI2, A1 => QI0, A2 => UQVN_N41, 
	A3 => EN, A4 => UQVN_N28);
UQVB_B45 : OR7
	PORT MAP (Z0 => UQVN_N39, A0 => HOLD2, A1 => LOAD2, A2 => UQVN_N38, 
	A3 => UQVN_N29, A4 => UQVN_N37, A5 => UQVN_N36, A6 => PS);
UQVB_B46 : AND7
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N45, A1 => QI1, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => EN, A5 => UQVN_N28, A6 => UQVN_N30);
UQVB_B47 : AND7
	PORT MAP (Z0 => UQVN_N29, A0 => QI3, A1 => QI1, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => EN, A5 => UQVN_N28, A6 => DNUP);
UQVB_B48 : AND4
	PORT MAP (Z0 => HOLD3, A0 => QI3, A1 => UQVN_N41, A2 => UQVN_N40, 
	A3 => UQVN_N28);
UQVB_B49 : AND7
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N44, A1 => UQVN_N43, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => EN, A5 => UQVN_N28, A6 => DNUP);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => CS);
UQVB_B51 : OR7
	PORT MAP (Z0 => UQVN_N34, A0 => HOLD3, A1 => LOAD3, A2 => UQVN_N33, 
	A3 => UQVN_N35, A4 => UQVN_N32, A5 => UQVN_N31, A6 => PS);
UQVB_B52 : AND7
	PORT MAP (Z0 => UQVN_N33, A0 => QI2, A1 => UQVN_N43, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => EN, A5 => UQVN_N28, A6 => UQVN_N30);
UQVB_B53 : AND5
	PORT MAP (Z0 => UQVN_N32, A0 => QI3, A1 => QI0, A2 => UQVN_N41, 
	A3 => EN, A4 => UQVN_N28);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => LD);
UQVB_B55 : AND5
	PORT MAP (Z0 => UQVN_N31, A0 => QI3, A1 => QI1, A2 => UQVN_N41, 
	A3 => EN, A4 => UQVN_N28);
UQVB_B56 : AND3
	PORT MAP (Z0 => LOAD3, A0 => D3, A1 => LD, A2 => UQVN_N28);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => QI3);
UQVB_B58 : FD21
	PORT MAP (Q0 => QI3, D0 => UQVN_N34, CLK => CLK, CD => CD);
UQVB_B59 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => DNUP);
UQVB_B60 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => QI2);
UQVB_B61 : FD21
	PORT MAP (Q0 => QI2, D0 => UQVN_N39, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for CMP2
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CMP2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        EQ : OUT std_logic
    );
END CMP2;


ARCHITECTURE lattice_arch OF CMP2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT NOR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR4 use  entity  lat_vhd.NOR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N8, A1 => B1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => UQVN_N6);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N7, A1 => B0);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => A0, A1 => UQVN_N5);
UQVB_B5 : NOR4
	PORT MAP (ZN0 => EQ, A0 => UQVN_N4, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => B0);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => B1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => A0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => A1);
END lattice_arch;
-- VHDL netlist for CMP4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CMP4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        EQ : OUT std_logic
    );
END CMP4;


ARCHITECTURE lattice_arch OF CMP4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT NOR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR8 use  entity  lat_vhd.NOR8(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => A2, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N15, A1 => B2);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => B2);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N16, A1 => B3);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => A2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => A3);
UQVB_B7 : NOR8
	PORT MAP (ZN0 => EQ, A0 => UQVN_N10, A1 => UQVN_N7, A2 => UQVN_N8, 
	A3 => UQVN_N9, A4 => UQVN_N3, A5 => UQVN_N4, A6 => UQVN_N5, 
	A7 => UQVN_N6);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N14, A1 => B1);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => A1, A1 => UQVN_N12);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N13, A1 => B0);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N10, A0 => A0, A1 => UQVN_N11);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => B0);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => B1);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => A0);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => A1);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => A3, A1 => UQVN_N2);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => B3);
END lattice_arch;
-- VHDL netlist for CMP8
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY CMP8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        EQ : OUT std_logic
    );
END CMP8;


ARCHITECTURE lattice_arch OF CMP8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT NOR16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR16 use  entity  lat_vhd.NOR16(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => A2, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N31, A1 => B2);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => B2);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N32, A1 => B3);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => A2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => A3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => A5, A1 => UQVN_N6);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => B5);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => A4, A1 => UQVN_N5);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N3, A1 => B4);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => B4);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N4, A1 => B5);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => A4);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => A5);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => A7);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => A6);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N9, A1 => B7);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => B6);
UQVB_B19 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N10, A1 => B6);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A6, A1 => UQVN_N8);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => B7);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => A7, A1 => UQVN_N7);
UQVB_B23 : NOR16
	PORT MAP (ZN0 => EQ, A0 => UQVN_N26, A1 => UQVN_N23, A2 => UQVN_N24, 
	A3 => UQVN_N25, A4 => UQVN_N22, A5 => UQVN_N21, A6 => UQVN_N15, 
	A7 => UQVN_N14, A8 => UQVN_N13, A9 => UQVN_N16, A10 => UQVN_N17, 
	A11 => UQVN_N18, A12 => UQVN_N11, A13 => UQVN_N12, A14 => UQVN_N20, 
	A15 => UQVN_N19);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N30, A1 => B1);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N24, A0 => A1, A1 => UQVN_N28);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N29, A1 => B0);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N26, A0 => A0, A1 => UQVN_N27);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => B0);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => B1);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => A0);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => A1);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => A3, A1 => UQVN_N2);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => B3);
END lattice_arch;
-- VHDL netlist for DEC2
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DEC2 IS 
    PORT (
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DEC2;


ARCHITECTURE lattice_arch OF DEC2 IS

  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => Z0, A0 => S0);
UQVB_B2 : BUF
	PORT MAP (Z0 => Z1, A0 => S0);
END lattice_arch;
-- VHDL netlist for DEC2E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DEC2E IS 
    PORT (
        EN : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DEC2E;


ARCHITECTURE lattice_arch OF DEC2E IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Z0, A0 => EN, A1 => UQVN_N1);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B3 : AND2
	PORT MAP (Z0 => Z1, A0 => EN, A1 => S0);
END lattice_arch;
-- VHDL netlist for DEC3
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DEC3 IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic
    );
END DEC3;


ARCHITECTURE lattice_arch OF DEC3 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N1);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S1);
UQVB_B3 : AND2
	PORT MAP (Z0 => Z1, A0 => S0, A1 => UQVN_N1);
UQVB_B4 : AND2
	PORT MAP (Z0 => Z2, A0 => UQVN_N2, A1 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
END lattice_arch;
-- VHDL netlist for DEC3E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DEC3E IS 
    PORT (
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic
    );
END DEC3E;


ARCHITECTURE lattice_arch OF DEC3E IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Z0, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N1);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z1, A0 => EN, A1 => S0, A2 => UQVN_N1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S1);
UQVB_B4 : AND3
	PORT MAP (Z0 => Z2, A0 => EN, A1 => UQVN_N2, A2 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
END lattice_arch;
-- VHDL netlist for DEC4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DEC4 IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DEC4;


ARCHITECTURE lattice_arch OF DEC4 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => Z3, A0 => S0, A1 => S1);
UQVB_B3 : AND2
	PORT MAP (Z0 => Z1, A0 => S0, A1 => UQVN_N1);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S1);
UQVB_B5 : AND2
	PORT MAP (Z0 => Z2, A0 => UQVN_N2, A1 => S1);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
END lattice_arch;
-- VHDL netlist for DEC4E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DEC4E IS 
    PORT (
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DEC4E;


ARCHITECTURE lattice_arch OF DEC4E IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Z0, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N1);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z3, A0 => EN, A1 => S0, A2 => S1);
UQVB_B3 : AND3
	PORT MAP (Z0 => Z1, A0 => EN, A1 => S0, A2 => UQVN_N1);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S1);
UQVB_B5 : AND3
	PORT MAP (Z0 => Z2, A0 => EN, A1 => UQVN_N2, A2 => S1);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX2
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX2 IS 
    PORT (
        A0 : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DMUX2;


ARCHITECTURE lattice_arch OF DMUX2 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => Z1, A0 => A0, A1 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX22
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX22 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        S0 : IN std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DMUX22;


ARCHITECTURE lattice_arch OF DMUX22 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Y0, A0 => A0, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B4 : AND2
	PORT MAP (Z0 => Y1, A0 => A1, A1 => UQVN_N2);
UQVB_B5 : AND2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX22E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX22E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DMUX22E;


ARCHITECTURE lattice_arch OF DMUX22E IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Y0, A0 => EN, A1 => A0, A2 => UQVN_N1);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B4 : AND3
	PORT MAP (Z0 => Y1, A0 => EN, A1 => A1, A2 => UQVN_N2);
UQVB_B5 : AND3
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A1, A2 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        W0 : OUT std_logic;
        W1 : OUT std_logic;
        X0 : OUT std_logic;
        X1 : OUT std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DMUX24;


ARCHITECTURE lattice_arch OF DMUX24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => W0, A0 => A0, A1 => UQVN_N1, A2 => UQVN_N2);
UQVB_B2 : AND3
	PORT MAP (Z0 => X0, A0 => A0, A1 => S0, A2 => UQVN_N2);
UQVB_B3 : AND3
	PORT MAP (Z0 => Y0, A0 => A0, A1 => UQVN_N1, A2 => S1);
UQVB_B4 : AND3
	PORT MAP (Z0 => Z0, A0 => A0, A1 => S0, A2 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
UQVB_B7 : AND3
	PORT MAP (Z0 => W1, A0 => A1, A1 => UQVN_N3, A2 => UQVN_N4);
UQVB_B8 : AND3
	PORT MAP (Z0 => X1, A0 => A1, A1 => S0, A2 => UQVN_N4);
UQVB_B9 : AND3
	PORT MAP (Z0 => Y1, A0 => A1, A1 => UQVN_N3, A2 => S1);
UQVB_B10 : AND3
	PORT MAP (Z0 => Z1, A0 => A1, A1 => S0, A2 => S1);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S1);
END lattice_arch;
-- VHDL netlist for DMUX24E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX24E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        W0 : OUT std_logic;
        W1 : OUT std_logic;
        X0 : OUT std_logic;
        X1 : OUT std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DMUX24E;


ARCHITECTURE lattice_arch OF DMUX24E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => W0, A0 => EN, A1 => A0, A2 => UQVN_N1, 
	A3 => UQVN_N2);
UQVB_B2 : AND4
	PORT MAP (Z0 => X0, A0 => EN, A1 => A0, A2 => S0, 
	A3 => UQVN_N2);
UQVB_B3 : AND4
	PORT MAP (Z0 => Y0, A0 => EN, A1 => A0, A2 => UQVN_N1, 
	A3 => S1);
UQVB_B4 : AND4
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => S0, 
	A3 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
UQVB_B7 : AND4
	PORT MAP (Z0 => W1, A0 => EN, A1 => A1, A2 => UQVN_N3, 
	A3 => UQVN_N4);
UQVB_B8 : AND4
	PORT MAP (Z0 => X1, A0 => EN, A1 => A1, A2 => S0, 
	A3 => UQVN_N4);
UQVB_B9 : AND4
	PORT MAP (Z0 => Y1, A0 => EN, A1 => A1, A2 => UQVN_N3, 
	A3 => S1);
UQVB_B10 : AND4
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A1, A2 => S0, 
	A3 => S1);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S1);
END lattice_arch;
-- VHDL netlist for DMUX2E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX2E IS 
    PORT (
        A0 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END DMUX2E;


ARCHITECTURE lattice_arch OF DMUX2E IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => UQVN_N1);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A0, A2 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX4 IS 
    PORT (
        A0 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DMUX4;


ARCHITECTURE lattice_arch OF DMUX4 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N1, A2 => UQVN_N2);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z1, A0 => A0, A1 => S0, A2 => UQVN_N2);
UQVB_B3 : AND3
	PORT MAP (Z0 => Z2, A0 => A0, A1 => UQVN_N1, A2 => S1);
UQVB_B4 : AND3
	PORT MAP (Z0 => Z3, A0 => A0, A1 => S0, A2 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
END lattice_arch;
-- VHDL netlist for DMUX42
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX42 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        S0 : IN std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Y2 : OUT std_logic;
        Y3 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DMUX42;


ARCHITECTURE lattice_arch OF DMUX42 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Y0, A0 => A0, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B4 : AND2
	PORT MAP (Z0 => Y1, A0 => A1, A1 => UQVN_N2);
UQVB_B5 : AND2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
UQVB_B7 : AND2
	PORT MAP (Z0 => Y3, A0 => A3, A1 => UQVN_N3);
UQVB_B8 : AND2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => S0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B10 : AND2
	PORT MAP (Z0 => Y2, A0 => A2, A1 => UQVN_N4);
UQVB_B11 : AND2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX42E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX42E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Y2 : OUT std_logic;
        Y3 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DMUX42E;


ARCHITECTURE lattice_arch OF DMUX42E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Y0, A0 => EN, A1 => A0, A2 => UQVN_N1);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B4 : AND3
	PORT MAP (Z0 => Y1, A0 => EN, A1 => A1, A2 => UQVN_N2);
UQVB_B5 : AND3
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A1, A2 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
UQVB_B7 : AND3
	PORT MAP (Z0 => Y3, A0 => EN, A1 => A3, A2 => UQVN_N3);
UQVB_B8 : AND3
	PORT MAP (Z0 => Z3, A0 => EN, A1 => A3, A2 => S0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B10 : AND3
	PORT MAP (Z0 => Y2, A0 => EN, A1 => A2, A2 => UQVN_N4);
UQVB_B11 : AND3
	PORT MAP (Z0 => Z2, A0 => EN, A1 => A2, A2 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX44
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        W0 : OUT std_logic;
        W1 : OUT std_logic;
        W2 : OUT std_logic;
        W3 : OUT std_logic;
        X0 : OUT std_logic;
        X1 : OUT std_logic;
        X2 : OUT std_logic;
        X3 : OUT std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Y2 : OUT std_logic;
        Y3 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DMUX44;


ARCHITECTURE lattice_arch OF DMUX44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => W0, A0 => A0, A1 => UQVN_N1, A2 => UQVN_N2);
UQVB_B2 : AND3
	PORT MAP (Z0 => X0, A0 => A0, A1 => S0, A2 => UQVN_N2);
UQVB_B3 : AND3
	PORT MAP (Z0 => Y0, A0 => A0, A1 => UQVN_N1, A2 => S1);
UQVB_B4 : AND3
	PORT MAP (Z0 => Z0, A0 => A0, A1 => S0, A2 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
UQVB_B7 : AND3
	PORT MAP (Z0 => W1, A0 => A1, A1 => UQVN_N3, A2 => UQVN_N4);
UQVB_B8 : AND3
	PORT MAP (Z0 => X1, A0 => A1, A1 => S0, A2 => UQVN_N4);
UQVB_B9 : AND3
	PORT MAP (Z0 => Y1, A0 => A1, A1 => UQVN_N3, A2 => S1);
UQVB_B10 : AND3
	PORT MAP (Z0 => Z1, A0 => A1, A1 => S0, A2 => S1);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S1);
UQVB_B13 : AND3
	PORT MAP (Z0 => W3, A0 => A3, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B14 : AND3
	PORT MAP (Z0 => X3, A0 => A3, A1 => S0, A2 => UQVN_N6);
UQVB_B15 : AND3
	PORT MAP (Z0 => Y3, A0 => A3, A1 => UQVN_N5, A2 => S1);
UQVB_B16 : AND3
	PORT MAP (Z0 => Z3, A0 => A3, A1 => S0, A2 => S1);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S1);
UQVB_B19 : AND3
	PORT MAP (Z0 => W2, A0 => A2, A1 => UQVN_N7, A2 => UQVN_N8);
UQVB_B20 : AND3
	PORT MAP (Z0 => X2, A0 => A2, A1 => S0, A2 => UQVN_N8);
UQVB_B21 : AND3
	PORT MAP (Z0 => Y2, A0 => A2, A1 => UQVN_N7, A2 => S1);
UQVB_B22 : AND3
	PORT MAP (Z0 => Z2, A0 => A2, A1 => S0, A2 => S1);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => S1);
END lattice_arch;
-- VHDL netlist for DMUX44E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX44E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        W0 : OUT std_logic;
        W1 : OUT std_logic;
        W2 : OUT std_logic;
        W3 : OUT std_logic;
        X0 : OUT std_logic;
        X1 : OUT std_logic;
        X2 : OUT std_logic;
        X3 : OUT std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Y2 : OUT std_logic;
        Y3 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DMUX44E;


ARCHITECTURE lattice_arch OF DMUX44E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => W0, A0 => EN, A1 => A0, A2 => UQVN_N1, 
	A3 => UQVN_N2);
UQVB_B2 : AND4
	PORT MAP (Z0 => X0, A0 => EN, A1 => A0, A2 => S0, 
	A3 => UQVN_N2);
UQVB_B3 : AND4
	PORT MAP (Z0 => Y0, A0 => EN, A1 => A0, A2 => UQVN_N1, 
	A3 => S1);
UQVB_B4 : AND4
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => S0, 
	A3 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
UQVB_B7 : AND4
	PORT MAP (Z0 => W1, A0 => EN, A1 => A1, A2 => UQVN_N3, 
	A3 => UQVN_N4);
UQVB_B8 : AND4
	PORT MAP (Z0 => X1, A0 => EN, A1 => A1, A2 => S0, 
	A3 => UQVN_N4);
UQVB_B9 : AND4
	PORT MAP (Z0 => Y1, A0 => EN, A1 => A1, A2 => UQVN_N3, 
	A3 => S1);
UQVB_B10 : AND4
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A1, A2 => S0, 
	A3 => S1);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S1);
UQVB_B13 : AND4
	PORT MAP (Z0 => W2, A0 => EN, A1 => A2, A2 => UQVN_N5, 
	A3 => UQVN_N6);
UQVB_B14 : AND4
	PORT MAP (Z0 => X2, A0 => EN, A1 => A2, A2 => S0, 
	A3 => UQVN_N6);
UQVB_B15 : AND4
	PORT MAP (Z0 => Y2, A0 => EN, A1 => A2, A2 => UQVN_N5, 
	A3 => S1);
UQVB_B16 : AND4
	PORT MAP (Z0 => Z2, A0 => EN, A1 => A2, A2 => S0, 
	A3 => S1);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S1);
UQVB_B19 : AND4
	PORT MAP (Z0 => W3, A0 => EN, A1 => A3, A2 => UQVN_N7, 
	A3 => UQVN_N8);
UQVB_B20 : AND4
	PORT MAP (Z0 => X3, A0 => EN, A1 => A3, A2 => S0, 
	A3 => UQVN_N8);
UQVB_B21 : AND4
	PORT MAP (Z0 => Y3, A0 => EN, A1 => A3, A2 => UQVN_N7, 
	A3 => S1);
UQVB_B22 : AND4
	PORT MAP (Z0 => Z3, A0 => EN, A1 => A3, A2 => S0, 
	A3 => S1);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => S1);
END lattice_arch;
-- VHDL netlist for DMUX4E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX4E IS 
    PORT (
        A0 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END DMUX4E;


ARCHITECTURE lattice_arch OF DMUX4E IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => UQVN_N1, 
	A3 => UQVN_N2);
UQVB_B2 : AND4
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A0, A2 => S0, 
	A3 => UQVN_N2);
UQVB_B3 : AND4
	PORT MAP (Z0 => Z2, A0 => EN, A1 => A0, A2 => UQVN_N1, 
	A3 => S1);
UQVB_B4 : AND4
	PORT MAP (Z0 => Z3, A0 => EN, A1 => A0, A2 => S0, 
	A3 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
END lattice_arch;
-- VHDL netlist for DMUX82
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX82 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        S0 : IN std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Y2 : OUT std_logic;
        Y3 : OUT std_logic;
        Y4 : OUT std_logic;
        Y5 : OUT std_logic;
        Y6 : OUT std_logic;
        Y7 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic
    );
END DMUX82;


ARCHITECTURE lattice_arch OF DMUX82 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Y0, A0 => A0, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B4 : AND2
	PORT MAP (Z0 => Y1, A0 => A1, A1 => UQVN_N2);
UQVB_B5 : AND2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
UQVB_B7 : AND2
	PORT MAP (Z0 => Y3, A0 => A3, A1 => UQVN_N3);
UQVB_B8 : AND2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => S0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B10 : AND2
	PORT MAP (Z0 => Y2, A0 => A2, A1 => UQVN_N4);
UQVB_B11 : AND2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B13 : AND2
	PORT MAP (Z0 => Y7, A0 => A7, A1 => UQVN_N5);
UQVB_B14 : AND2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => S0);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B16 : AND2
	PORT MAP (Z0 => Y6, A0 => A6, A1 => UQVN_N6);
UQVB_B17 : AND2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => S0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S0);
UQVB_B19 : AND2
	PORT MAP (Z0 => Y4, A0 => A4, A1 => UQVN_N7);
UQVB_B20 : AND2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => S0);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B22 : AND2
	PORT MAP (Z0 => Y5, A0 => A5, A1 => UQVN_N8);
UQVB_B23 : AND2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => S0);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => S0);
END lattice_arch;
-- VHDL netlist for DMUX82E
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY DMUX82E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Y0 : OUT std_logic;
        Y1 : OUT std_logic;
        Y2 : OUT std_logic;
        Y3 : OUT std_logic;
        Y4 : OUT std_logic;
        Y5 : OUT std_logic;
        Y6 : OUT std_logic;
        Y7 : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic
    );
END DMUX82E;


ARCHITECTURE lattice_arch OF DMUX82E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => Y0, A0 => EN, A1 => A0, A2 => UQVN_N1);
UQVB_B2 : AND3
	PORT MAP (Z0 => Z0, A0 => EN, A1 => A0, A2 => S0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B4 : AND3
	PORT MAP (Z0 => Y1, A0 => EN, A1 => A1, A2 => UQVN_N2);
UQVB_B5 : AND3
	PORT MAP (Z0 => Z1, A0 => EN, A1 => A1, A2 => S0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S0);
UQVB_B7 : AND3
	PORT MAP (Z0 => Y3, A0 => EN, A1 => A3, A2 => UQVN_N3);
UQVB_B8 : AND3
	PORT MAP (Z0 => Z3, A0 => EN, A1 => A3, A2 => S0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S0);
UQVB_B10 : AND3
	PORT MAP (Z0 => Y2, A0 => EN, A1 => A2, A2 => UQVN_N4);
UQVB_B11 : AND3
	PORT MAP (Z0 => Z2, A0 => EN, A1 => A2, A2 => S0);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B13 : AND3
	PORT MAP (Z0 => Y7, A0 => EN, A1 => A7, A2 => UQVN_N5);
UQVB_B14 : AND3
	PORT MAP (Z0 => Z7, A0 => EN, A1 => A7, A2 => S0);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B16 : AND3
	PORT MAP (Z0 => Y6, A0 => EN, A1 => A6, A2 => UQVN_N6);
UQVB_B17 : AND3
	PORT MAP (Z0 => Z6, A0 => EN, A1 => A6, A2 => S0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S0);
UQVB_B19 : AND3
	PORT MAP (Z0 => Y4, A0 => EN, A1 => A4, A2 => UQVN_N7);
UQVB_B20 : AND3
	PORT MAP (Z0 => Z4, A0 => EN, A1 => A4, A2 => S0);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B22 : AND3
	PORT MAP (Z0 => Y5, A0 => EN, A1 => A5, A2 => UQVN_N8);
UQVB_B23 : AND3
	PORT MAP (Z0 => Z5, A0 => EN, A1 => A5, A2 => S0);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => S0);
END lattice_arch;
-- VHDL netlist for F3ADD
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY F3ADD IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        G012 : OUT std_logic;
        P012 : OUT std_logic
    );
END F3ADD;


ARCHITECTURE lattice_arch OF F3ADD IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => CI);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B2);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => A0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N40, A1 => CI);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => UQVN_N43);
UQVB_B7 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N3);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N37, A1 => B1, A2 => UQVN_N40);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N41, A1 => B0, A2 => CI);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => A0, A1 => UQVN_N41, A2 => CI);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B1, A1 => UQVN_N40, A2 => UQVN_N43);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N37, A1 => B1, A2 => UQVN_N43);
UQVB_B14 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N8);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => UQVN_N41, A2 => B0);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => A0, A1 => A1, A2 => A2, 
	A3 => B0);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A1, A1 => A2, A2 => B1);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => A0, A1 => A2, A2 => B0, 
	A3 => B1);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A2, A1 => B2);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B2);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => A1, A1 => B1, A2 => B2);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => A0, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B24 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16, A6 => UQVN_N17);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N37, A1 => UQVN_N40);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N38, A1 => UQVN_N41);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N39, A1 => UQVN_N42);
UQVB_B28 : NOR3
	PORT MAP (ZN0 => P012, A0 => UQVN_N20, A1 => UQVN_N18, A2 => UQVN_N19);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => B0);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A1);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A2);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N34);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N41, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N38, A1 => UQVN_N40, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N37, A1 => UQVN_N38, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => B0, A1 => B1, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => A0, A1 => B1, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A1, A1 => B0, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => A0, A1 => A1, A2 => UQVN_N42, 
	A3 => CI);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => A0, A1 => B0, A2 => B1, 
	A3 => UQVN_N42);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => A1, A1 => B1, A2 => UQVN_N42);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => A0, A1 => A1, A2 => B0, 
	A3 => UQVN_N42);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N37, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => B2);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N38, A1 => UQVN_N41, A2 => B2);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N37, A1 => UQVN_N38, A2 => UQVN_N40, 
	A3 => B2);
UQVB_B47 : OR12
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N28, A5 => UQVN_N27, A6 => UQVN_N26, 
	A7 => UQVN_N25, A8 => UQVN_N24, A9 => UQVN_N23, A10 => UQVN_N22, 
	A11 => UQVN_N21);
UQVB_B48 : OR3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N33, A1 => UQVN_N35, A2 => UQVN_N36);
END lattice_arch;
-- VHDL netlist for F3SUB
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY F3SUB IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        BI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        G012 : OUT std_logic;
        P012 : OUT std_logic
    );
END F3SUB;


ARCHITECTURE lattice_arch OF F3SUB IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => BI);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B2);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => A0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N40, A1 => BI);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => UQVN_N43);
UQVB_B7 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B8 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N3);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => A0, A1 => B1, A2 => UQVN_N40);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N41, A1 => B0, A2 => BI);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N37, A1 => UQVN_N41, A2 => BI);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B1, A1 => UQVN_N40, A2 => UQVN_N43);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A0, A1 => B1, A2 => UQVN_N43);
UQVB_B14 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N8);
UQVB_B15 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N10);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N37, A1 => UQVN_N41, A2 => B0);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N37, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N38, A1 => B1, A2 => B2);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N37, A1 => UQVN_N39, A2 => B0, 
	A3 => B1);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N39, A1 => B2);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N37, A1 => UQVN_N38, A2 => B0, 
	A3 => B2);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N38, A1 => UQVN_N39, A2 => B1);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N37, A1 => UQVN_N38, A2 => UQVN_N39, 
	A3 => B0);
UQVB_B24 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N15, A5 => UQVN_N16, A6 => UQVN_N17);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => A0, A1 => UQVN_N40);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => A1, A1 => UQVN_N41);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => A2, A1 => UQVN_N42);
UQVB_B28 : NOR3
	PORT MAP (ZN0 => P012, A0 => UQVN_N20, A1 => UQVN_N18, A2 => UQVN_N19);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => B0);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A1);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A2);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N34);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => A0, A1 => A1, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N37, A1 => UQVN_N38, A2 => UQVN_N42, 
	A3 => BI);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => A0, A1 => A1, A2 => UQVN_N40, 
	A3 => B2);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => A1, A1 => UQVN_N40, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N37, A1 => UQVN_N38, A2 => B0, 
	A3 => UQVN_N42);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N38, A1 => B0, A2 => UQVN_N42, 
	A3 => BI);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A0, A1 => UQVN_N41, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => A0, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => B2);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B2, 
	A3 => UQVN_N43);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N38, A1 => UQVN_N42, A2 => B1);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N37, A1 => B1, A2 => UQVN_N42, 
	A3 => BI);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N37, A1 => B0, A2 => B1, 
	A3 => UQVN_N42);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => A1, A1 => UQVN_N41, A2 => B2);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => B0, A1 => B1, A2 => UQVN_N42, 
	A3 => BI);
UQVB_B47 : OR12
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N28, A5 => UQVN_N27, A6 => UQVN_N26, 
	A7 => UQVN_N25, A8 => UQVN_N24, A9 => UQVN_N23, A10 => UQVN_N22, 
	A11 => UQVN_N21);
UQVB_B48 : OR3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N33, A1 => UQVN_N35, A2 => UQVN_N36);
END lattice_arch;
-- VHDL netlist for FD14
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD14;


ARCHITECTURE lattice_arch OF FD14 IS

  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q3, D0 => D3, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => Q2, D0 => D2, CLK => CLK);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q1, D0 => D1, CLK => CLK);
UQVB_B4 : FD11
	PORT MAP (Q0 => Q0, D0 => D0, CLK => CLK);
END lattice_arch;
-- VHDL netlist for FD18
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD18 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD18;


ARCHITECTURE lattice_arch OF FD18 IS

  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q3, D0 => D3, CLK => CLK);
UQVB_B2 : FD11
	PORT MAP (Q0 => Q2, D0 => D2, CLK => CLK);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q1, D0 => D1, CLK => CLK);
UQVB_B4 : FD11
	PORT MAP (Q0 => Q0, D0 => D0, CLK => CLK);
UQVB_B5 : FD11
	PORT MAP (Q0 => Q4, D0 => D4, CLK => CLK);
UQVB_B6 : FD11
	PORT MAP (Q0 => Q5, D0 => D5, CLK => CLK);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q6, D0 => D6, CLK => CLK);
UQVB_B8 : FD11
	PORT MAP (Q0 => Q7, D0 => D7, CLK => CLK);
END lattice_arch;
-- VHDL netlist for FD24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD24 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD24;


ARCHITECTURE lattice_arch OF FD24 IS

  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => Q3, D0 => D3, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => Q2, D0 => D2, CLK => CLK, CD => CD);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q1, D0 => D1, CLK => CLK, CD => CD);
UQVB_B4 : FD21
	PORT MAP (Q0 => Q0, D0 => D0, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for FD28
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD28 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD28;


ARCHITECTURE lattice_arch OF FD28 IS

  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => Q3, D0 => D3, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => Q2, D0 => D2, CLK => CLK, CD => CD);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q1, D0 => D1, CLK => CLK, CD => CD);
UQVB_B4 : FD21
	PORT MAP (Q0 => Q0, D0 => D0, CLK => CLK, CD => CD);
UQVB_B5 : FD21
	PORT MAP (Q0 => Q6, D0 => D6, CLK => CLK, CD => CD);
UQVB_B6 : FD21
	PORT MAP (Q0 => Q5, D0 => D5, CLK => CLK, CD => CD);
UQVB_B7 : FD21
	PORT MAP (Q0 => Q4, D0 => D4, CLK => CLK, CD => CD);
UQVB_B8 : FD21
	PORT MAP (Q0 => Q7, D0 => D7, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for FD31
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD31 IS 
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        Q0 : OUT std_logic
    );
END FD31;


ARCHITECTURE lattice_arch OF FD31 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => D0, A1 => PS);
END lattice_arch;
-- VHDL netlist for FD34
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD34;


ARCHITECTURE lattice_arch OF FD34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => PS);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => D2, A1 => PS);
UQVB_B5 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, CLK => CLK);
UQVB_B6 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => PS);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, CLK => CLK);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => PS);
END lattice_arch;
-- VHDL netlist for FD38
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD38;


ARCHITECTURE lattice_arch OF FD38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q7, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => D7, A1 => PS);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q6, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => D6, A1 => PS);
UQVB_B5 : FD11
	PORT MAP (Q0 => Q5, D0 => UQVN_N3, CLK => CLK);
UQVB_B6 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => D5, A1 => PS);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q4, D0 => UQVN_N4, CLK => CLK);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => D4, A1 => PS);
UQVB_B9 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, CLK => CLK);
UQVB_B10 : OR2
	PORT MAP (Z0 => UQVN_N5, A0 => D2, A1 => PS);
UQVB_B11 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N6, CLK => CLK);
UQVB_B12 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => D3, A1 => PS);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N7, CLK => CLK);
UQVB_B14 : OR2
	PORT MAP (Z0 => UQVN_N7, A0 => D1, A1 => PS);
UQVB_B15 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N8, CLK => CLK);
UQVB_B16 : OR2
	PORT MAP (Z0 => UQVN_N8, A0 => D0, A1 => PS);
END lattice_arch;
-- VHDL netlist for FD41
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD41 IS 
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END FD41;


ARCHITECTURE lattice_arch OF FD41 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => D0, A1 => PS);
END lattice_arch;
-- VHDL netlist for FD44
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD44;


ARCHITECTURE lattice_arch OF FD44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => PS);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => D2, A1 => PS);
UQVB_B5 : FD21
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B6 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => PS);
UQVB_B7 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => PS);
END lattice_arch;
-- VHDL netlist for FD48
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD48;


ARCHITECTURE lattice_arch OF FD48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => PS);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => D2, A1 => PS);
UQVB_B5 : FD21
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B6 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => D1, A1 => PS);
UQVB_B7 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => PS);
UQVB_B9 : FD21
	PORT MAP (Q0 => Q7, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B10 : OR2
	PORT MAP (Z0 => UQVN_N5, A0 => D7, A1 => PS);
UQVB_B11 : FD21
	PORT MAP (Q0 => Q6, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B12 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => D6, A1 => PS);
UQVB_B13 : FD21
	PORT MAP (Q0 => Q5, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B14 : OR2
	PORT MAP (Z0 => UQVN_N7, A0 => D5, A1 => PS);
UQVB_B15 : FD21
	PORT MAP (Q0 => Q4, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B16 : OR2
	PORT MAP (Z0 => UQVN_N8, A0 => D4, A1 => PS);
END lattice_arch;
-- VHDL netlist for FD51
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD51 IS 
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic
    );
END FD51;


ARCHITECTURE lattice_arch OF FD51 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N1, A1 => PS);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => CS);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => D0, A1 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for FD54
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD54 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD54;


ARCHITECTURE lattice_arch OF FD54 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N1, A1 => PS);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => CS);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => UQVN_N3);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N4, A1 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => CS);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, CLK => CLK);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => D2, A1 => UQVN_N6);
UQVB_B9 : OR2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N7, A1 => PS);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => CS);
UQVB_B11 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N8, CLK => CLK);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => D1, A1 => UQVN_N9);
UQVB_B13 : OR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N10, A1 => PS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CS);
UQVB_B15 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N11, CLK => CLK);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N10, A0 => D0, A1 => UQVN_N12);
END lattice_arch;
-- VHDL netlist for FD58
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD58 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD58;


ARCHITECTURE lattice_arch OF FD58 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N1, A1 => PS);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => CS);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => UQVN_N3);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N4, A1 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => CS);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N5, CLK => CLK);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => D2, A1 => UQVN_N6);
UQVB_B9 : OR2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N7, A1 => PS);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => CS);
UQVB_B11 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N8, CLK => CLK);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => D1, A1 => UQVN_N9);
UQVB_B13 : OR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N10, A1 => PS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CS);
UQVB_B15 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N11, CLK => CLK);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N10, A0 => D0, A1 => UQVN_N12);
UQVB_B17 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N13, A1 => PS);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => CS);
UQVB_B19 : FD11
	PORT MAP (Q0 => Q7, D0 => UQVN_N14, CLK => CLK);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => D7, A1 => UQVN_N15);
UQVB_B21 : OR2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N16, A1 => PS);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => CS);
UQVB_B23 : FD11
	PORT MAP (Q0 => Q6, D0 => UQVN_N17, CLK => CLK);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => D6, A1 => UQVN_N18);
UQVB_B25 : OR2
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N19, A1 => PS);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => CS);
UQVB_B27 : FD11
	PORT MAP (Q0 => Q5, D0 => UQVN_N20, CLK => CLK);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D5, A1 => UQVN_N21);
UQVB_B29 : OR2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N22, A1 => PS);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => CS);
UQVB_B31 : FD11
	PORT MAP (Q0 => Q4, D0 => UQVN_N23, CLK => CLK);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => D4, A1 => UQVN_N24);
END lattice_arch;
-- VHDL netlist for FD61
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD61 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FD61;


ARCHITECTURE lattice_arch OF FD61 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI0, A1 => TE);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for FD64
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD64 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        CLK : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD64;


ARCHITECTURE lattice_arch OF FD64 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TE);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D2);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI2, A1 => TE);
UQVB_B8 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => CLK);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15);
END lattice_arch;
-- VHDL netlist for FD68
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD68 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        CLK : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD68;


ARCHITECTURE lattice_arch OF FD68 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TE);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D2);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI2, A1 => TE);
UQVB_B8 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => CLK);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N17, A1 => D6);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => TI6, A1 => TE);
UQVB_B23 : FD11
	PORT MAP (Q0 => Q6, D0 => UQVN_N18, CLK => CLK);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TE);
UQVB_B25 : OR2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N21, A1 => D5);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N24, A0 => TI5, A1 => TE);
UQVB_B28 : FD11
	PORT MAP (Q0 => Q5, D0 => UQVN_N22, CLK => CLK);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => TE);
UQVB_B30 : OR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N24, A1 => UQVN_N23);
UQVB_B31 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N25, A1 => D4);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => TI4, A1 => TE);
UQVB_B33 : FD11
	PORT MAP (Q0 => Q4, D0 => UQVN_N26, CLK => CLK);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => TE);
UQVB_B35 : OR2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N28, A1 => UQVN_N27);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N29, A1 => D7);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => TI7, A1 => TE);
UQVB_B38 : FD11
	PORT MAP (Q0 => Q7, D0 => UQVN_N30, CLK => CLK);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => TE);
UQVB_B40 : OR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N31);
END lattice_arch;
-- VHDL netlist for FD71
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD71 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FD71;


ARCHITECTURE lattice_arch OF FD71 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI0, A1 => TE);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for FD74
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD74 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD74;


ARCHITECTURE lattice_arch OF FD74 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TE);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D2);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI2, A1 => TE);
UQVB_B8 : FD21
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD21
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15);
END lattice_arch;
-- VHDL netlist for FD78
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD78 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD78;


ARCHITECTURE lattice_arch OF FD78 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TE);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D2);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI2, A1 => TE);
UQVB_B8 : FD21
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD21
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR2
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N17, A1 => D6);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => TI6, A1 => TE);
UQVB_B23 : FD21
	PORT MAP (Q0 => Q6, D0 => UQVN_N18, CLK => CLK, CD => CD);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TE);
UQVB_B25 : OR2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N21, A1 => D5);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N24, A0 => TI5, A1 => TE);
UQVB_B28 : FD21
	PORT MAP (Q0 => Q5, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => TE);
UQVB_B30 : OR2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N24, A1 => UQVN_N23);
UQVB_B31 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N25, A1 => D4);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => TI4, A1 => TE);
UQVB_B33 : FD21
	PORT MAP (Q0 => Q4, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => TE);
UQVB_B35 : OR2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N28, A1 => UQVN_N27);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N29, A1 => D7);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => TI7, A1 => TE);
UQVB_B38 : FD21
	PORT MAP (Q0 => Q7, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => TE);
UQVB_B40 : OR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N31);
END lattice_arch;
-- VHDL netlist for FD81
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD81 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FD81;


ARCHITECTURE lattice_arch OF FD81 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI0, A1 => TE);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3, A2 => PS);
END lattice_arch;
-- VHDL netlist for FD84
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD84 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD84;


ARCHITECTURE lattice_arch OF FD84 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D2);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI2, A1 => TE);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3, A2 => PS);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI3, A1 => TE);
UQVB_B8 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N6, CLK => CLK);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7, A2 => PS);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11, A2 => PS);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15, A2 => PS);
END lattice_arch;
-- VHDL netlist for FD88
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD88 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD88;


ARCHITECTURE lattice_arch OF FD88 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D7);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI7, A1 => TE);
UQVB_B3 : FD11
	PORT MAP (Q0 => Q7, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3, A2 => PS);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D6);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI6, A1 => TE);
UQVB_B8 : FD11
	PORT MAP (Q0 => Q6, D0 => UQVN_N6, CLK => CLK);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7, A2 => PS);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D5);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI5, A1 => TE);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q5, D0 => UQVN_N10, CLK => CLK);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11, A2 => PS);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D4);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI4, A1 => TE);
UQVB_B18 : FD11
	PORT MAP (Q0 => Q4, D0 => UQVN_N14, CLK => CLK);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15, A2 => PS);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N17, A1 => D2);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => TI2, A1 => TE);
UQVB_B23 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N18, CLK => CLK);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TE);
UQVB_B25 : OR3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19, A2 => PS);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N21, A1 => D3);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N24, A0 => TI3, A1 => TE);
UQVB_B28 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N22, CLK => CLK);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => TE);
UQVB_B30 : OR3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N24, A1 => UQVN_N23, A2 => PS);
UQVB_B31 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N25, A1 => D1);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => TI1, A1 => TE);
UQVB_B33 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N26, CLK => CLK);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => TE);
UQVB_B35 : OR3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N28, A1 => UQVN_N27, A2 => PS);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N29, A1 => D0);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => TI0, A1 => TE);
UQVB_B38 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N30, CLK => CLK);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => TE);
UQVB_B40 : OR3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N31, A2 => PS);
END lattice_arch;
-- VHDL netlist for FD91
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD91 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FD91;


ARCHITECTURE lattice_arch OF FD91 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI0, A1 => TE);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3, A2 => PS);
END lattice_arch;
-- VHDL netlist for FD94
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD94 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FD94;


ARCHITECTURE lattice_arch OF FD94 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TE);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3, A2 => PS);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D2);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI2, A1 => TE);
UQVB_B8 : FD21
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7, A2 => PS);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD21
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11, A2 => PS);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15, A2 => PS);
END lattice_arch;
-- VHDL netlist for FD98
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FD98 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FD98;


ARCHITECTURE lattice_arch OF FD98 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N1, A1 => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TE);
UQVB_B3 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B5 : OR3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N3, A2 => PS);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N5, A1 => D2);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => TI2, A1 => TE);
UQVB_B8 : FD21
	PORT MAP (Q0 => Q2, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => TE);
UQVB_B10 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N7, A2 => PS);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N9, A1 => D1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI1, A1 => TE);
UQVB_B13 : FD21
	PORT MAP (Q0 => Q1, D0 => UQVN_N10, CLK => CLK, CD => CD);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TE);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N12, A1 => UQVN_N11, A2 => PS);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N13, A1 => D0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => TI0, A1 => TE);
UQVB_B18 : FD21
	PORT MAP (Q0 => Q0, D0 => UQVN_N14, CLK => CLK, CD => CD);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => TE);
UQVB_B20 : OR3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N15, A2 => PS);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N17, A1 => D7);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => TI7, A1 => TE);
UQVB_B23 : FD21
	PORT MAP (Q0 => Q7, D0 => UQVN_N18, CLK => CLK, CD => CD);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TE);
UQVB_B25 : OR3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19, A2 => PS);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N21, A1 => D6);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N24, A0 => TI6, A1 => TE);
UQVB_B28 : FD21
	PORT MAP (Q0 => Q6, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => TE);
UQVB_B30 : OR3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N24, A1 => UQVN_N23, A2 => PS);
UQVB_B31 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N25, A1 => D5);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => TI5, A1 => TE);
UQVB_B33 : FD21
	PORT MAP (Q0 => Q5, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => TE);
UQVB_B35 : OR3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N28, A1 => UQVN_N27, A2 => PS);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N29, A1 => D4);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => TI4, A1 => TE);
UQVB_B38 : FD21
	PORT MAP (Q0 => Q4, D0 => UQVN_N30, CLK => CLK, CD => CD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => TE);
UQVB_B40 : OR3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N31, A2 => PS);
END lattice_arch;
-- VHDL netlist for FDA1
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FDA1 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FDA1;


ARCHITECTURE lattice_arch OF FDA1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N3, CLK => CLK);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N4, A2 => PS);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N1, A1 => D0, A2 => UQVN_N2);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => TI0, A1 => TE, A2 => UQVN_N2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CS);
END lattice_arch;
-- VHDL netlist for FDA4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FDA4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FDA4;


ARCHITECTURE lattice_arch OF FDA4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, CLK => CLK);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N4, A2 => PS);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N1, A1 => D3, A2 => UQVN_N2);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => TI3, A1 => TE, A2 => UQVN_N2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CS);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N8, CLK => CLK);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => TE);
UQVB_B9 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N9, A2 => PS);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N6, A1 => D2, A2 => UQVN_N7);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => TI2, A1 => TE, A2 => UQVN_N7);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => CS);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N13, CLK => CLK);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => TE);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N15, A1 => UQVN_N14, A2 => PS);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N11, A1 => D1, A2 => UQVN_N12);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => TI1, A1 => TE, A2 => UQVN_N12);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CS);
UQVB_B19 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N18, CLK => CLK);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => TE);
UQVB_B21 : OR3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19, A2 => PS);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N16, A1 => D0, A2 => UQVN_N17);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => TI0, A1 => TE, A2 => UQVN_N17);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => CS);
END lattice_arch;
-- VHDL netlist for FDA8
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FDA8 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FDA8;


ARCHITECTURE lattice_arch OF FDA8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, CLK => CLK);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N4, A2 => PS);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N1, A1 => D3, A2 => UQVN_N2);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => TI3, A1 => TE, A2 => UQVN_N2);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CS);
UQVB_B7 : FD11
	PORT MAP (Q0 => Q2, D0 => UQVN_N8, CLK => CLK);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => TE);
UQVB_B9 : OR3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N9, A2 => PS);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N6, A1 => D2, A2 => UQVN_N7);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => TI2, A1 => TE, A2 => UQVN_N7);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => CS);
UQVB_B13 : FD11
	PORT MAP (Q0 => Q1, D0 => UQVN_N13, CLK => CLK);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => TE);
UQVB_B15 : OR3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N15, A1 => UQVN_N14, A2 => PS);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N11, A1 => D1, A2 => UQVN_N12);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => TI1, A1 => TE, A2 => UQVN_N12);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CS);
UQVB_B19 : FD11
	PORT MAP (Q0 => Q0, D0 => UQVN_N18, CLK => CLK);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => TE);
UQVB_B21 : OR3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19, A2 => PS);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N16, A1 => D0, A2 => UQVN_N17);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => TI0, A1 => TE, A2 => UQVN_N17);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => CS);
UQVB_B25 : FD11
	PORT MAP (Q0 => Q7, D0 => UQVN_N23, CLK => CLK);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => TE);
UQVB_B27 : OR3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N25, A1 => UQVN_N24, A2 => PS);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N21, A1 => D7, A2 => UQVN_N22);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => TI7, A1 => TE, A2 => UQVN_N22);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CS);
UQVB_B31 : FD11
	PORT MAP (Q0 => Q6, D0 => UQVN_N28, CLK => CLK);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => TE);
UQVB_B33 : OR3
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N30, A1 => UQVN_N29, A2 => PS);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N26, A1 => D6, A2 => UQVN_N27);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => TI6, A1 => TE, A2 => UQVN_N27);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => CS);
UQVB_B37 : FD11
	PORT MAP (Q0 => Q5, D0 => UQVN_N33, CLK => CLK);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => TE);
UQVB_B39 : OR3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N35, A1 => UQVN_N34, A2 => PS);
UQVB_B40 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N31, A1 => D5, A2 => UQVN_N32);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => TI5, A1 => TE, A2 => UQVN_N32);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => CS);
UQVB_B43 : FD11
	PORT MAP (Q0 => Q4, D0 => UQVN_N38, CLK => CLK);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => TE);
UQVB_B45 : OR3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N39, A2 => PS);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N36, A1 => D4, A2 => UQVN_N37);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N40, A0 => TI4, A1 => TE, A2 => UQVN_N37);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => CS);
END lattice_arch;
-- VHDL netlist for FDB1
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FDB1 IS 
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        SD : IN std_logic;
        Q0 : OUT std_logic
    );
END FDB1;


ARCHITECTURE lattice_arch OF FDB1 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N1, CLK => CLK, CD => SD);
UQVB_B2 : INV
	PORT MAP (ZN0 => Q0, A0 => UQVN_N2);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => D0);
END lattice_arch;
-- VHDL netlist for FDB4
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FDB4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CLK : IN std_logic;
        SD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END FDB4;


ARCHITECTURE lattice_arch OF FDB4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N1, CLK => CLK, CD => SD);
UQVB_B2 : INV
	PORT MAP (ZN0 => Q3, A0 => UQVN_N2);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => D3);
UQVB_B4 : FD21
	PORT MAP (Q0 => UQVN_N4, D0 => UQVN_N3, CLK => CLK, CD => SD);
UQVB_B5 : INV
	PORT MAP (ZN0 => Q2, A0 => UQVN_N4);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => D2);
UQVB_B7 : FD21
	PORT MAP (Q0 => UQVN_N6, D0 => UQVN_N5, CLK => CLK, CD => SD);
UQVB_B8 : INV
	PORT MAP (ZN0 => Q1, A0 => UQVN_N6);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => D1);
UQVB_B10 : FD21
	PORT MAP (Q0 => UQVN_N8, D0 => UQVN_N7, CLK => CLK, CD => SD);
UQVB_B11 : INV
	PORT MAP (ZN0 => Q0, A0 => UQVN_N8);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => D0);
END lattice_arch;
-- VHDL netlist for FDB8
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FDB8 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CLK : IN std_logic;
        SD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END FDB8;


ARCHITECTURE lattice_arch OF FDB8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N1, CLK => CLK, CD => SD);
UQVB_B2 : INV
	PORT MAP (ZN0 => Q3, A0 => UQVN_N2);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => D3);
UQVB_B4 : FD21
	PORT MAP (Q0 => UQVN_N4, D0 => UQVN_N3, CLK => CLK, CD => SD);
UQVB_B5 : INV
	PORT MAP (ZN0 => Q2, A0 => UQVN_N4);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => D2);
UQVB_B7 : FD21
	PORT MAP (Q0 => UQVN_N6, D0 => UQVN_N5, CLK => CLK, CD => SD);
UQVB_B8 : INV
	PORT MAP (ZN0 => Q1, A0 => UQVN_N6);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => D1);
UQVB_B10 : FD21
	PORT MAP (Q0 => UQVN_N8, D0 => UQVN_N7, CLK => CLK, CD => SD);
UQVB_B11 : INV
	PORT MAP (ZN0 => Q0, A0 => UQVN_N8);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => D0);
UQVB_B13 : FD21
	PORT MAP (Q0 => UQVN_N10, D0 => UQVN_N9, CLK => CLK, CD => SD);
UQVB_B14 : INV
	PORT MAP (ZN0 => Q6, A0 => UQVN_N10);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => D6);
UQVB_B16 : FD21
	PORT MAP (Q0 => UQVN_N12, D0 => UQVN_N11, CLK => CLK, CD => SD);
UQVB_B17 : INV
	PORT MAP (ZN0 => Q5, A0 => UQVN_N12);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => D5);
UQVB_B19 : FD21
	PORT MAP (Q0 => UQVN_N14, D0 => UQVN_N13, CLK => CLK, CD => SD);
UQVB_B20 : INV
	PORT MAP (ZN0 => Q4, A0 => UQVN_N14);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => D4);
UQVB_B22 : FD21
	PORT MAP (Q0 => UQVN_N16, D0 => UQVN_N15, CLK => CLK, CD => SD);
UQVB_B23 : INV
	PORT MAP (ZN0 => Q7, A0 => UQVN_N16);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => D7);
END lattice_arch;
-- VHDL netlist for FJK11
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FJK11 IS 
    PORT (
        J0 : IN std_logic;
        K0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
END FJK11;


ARCHITECTURE lattice_arch OF FJK11 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N4, CLK => CLK);
UQVB_B2 : NAND2
	PORT MAP (ZN0 => UQVN_N1, A0 => UQVN_N3, A1 => J0);
UQVB_B3 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N3, A1 => K0);
UQVB_B4 : NAND2
	PORT MAP (ZN0 => UQVN_N4, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => UQVN_N5);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
END lattice_arch;
-- VHDL netlist for FJK21
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FJK21 IS 
    PORT (
        J0 : IN std_logic;
        K0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END FJK21;


ARCHITECTURE lattice_arch OF FJK21 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N4, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B2 : NAND2
	PORT MAP (ZN0 => UQVN_N1, A0 => UQVN_N3, A1 => J0);
UQVB_B3 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N3, A1 => K0);
UQVB_B4 : NAND2
	PORT MAP (ZN0 => UQVN_N5, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => UQVN_N4);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N4);
END lattice_arch;
-- VHDL netlist for FJK31
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FJK31 IS 
    PORT (
        J0 : IN std_logic;
        K0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FJK31;


ARCHITECTURE lattice_arch OF FJK31 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B2 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
UQVB_B3 : FD11
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N7, CLK => CLK);
UQVB_B4 : NAND2
	PORT MAP (ZN0 => UQVN_N2, A0 => UQVN_N4, A1 => J0);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N4, A1 => K0);
UQVB_B6 : NAND2
	PORT MAP (ZN0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => UQVN_N5);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => TI0, A1 => TE);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for FJK41
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FJK41 IS 
    PORT (
        J0 : IN std_logic;
        K0 : IN std_logic;
        TI0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        TE : IN std_logic;
        Q0 : OUT std_logic
    );
END FJK41;


ARCHITECTURE lattice_arch OF FJK41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => TE);
UQVB_B2 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
UQVB_B3 : FD21
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B4 : NAND2
	PORT MAP (ZN0 => UQVN_N2, A0 => UQVN_N4, A1 => J0);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N4, A1 => K0);
UQVB_B6 : NAND2
	PORT MAP (ZN0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => UQVN_N5);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => TI0, A1 => TE);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N6, A1 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for FJK51
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FJK51 IS 
    PORT (
        J0 : IN std_logic;
        K0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END FJK51;


ARCHITECTURE lattice_arch OF FJK51 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B2 : NAND2
	PORT MAP (ZN0 => UQVN_N5, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B3 : NAND2
	PORT MAP (ZN0 => UQVN_N1, A0 => UQVN_N4, A1 => J0);
UQVB_B4 : OR2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N4, A1 => K0);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => UQVN_N3);
UQVB_B6 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N5, A1 => PS);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for FT11
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FT11 IS 
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END FT11;


ARCHITECTURE lattice_arch OF FT11 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
UQVB_B3 : XOR2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => D0);
END lattice_arch;
-- VHDL netlist for FT21
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY FT21 IS 
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic
    );
END FT21;


ARCHITECTURE lattice_arch OF FT21 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N3, CLK => CLK);
UQVB_B2 : XOR2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => D0);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => CS);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N5, A1 => UQVN_N1);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
UQVB_B6 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N4, A1 => PS);
END lattice_arch;
-- VHDL netlist for IB11
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IB11 IS 
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
END IB11;


ARCHITECTURE lattice_arch OF IB11 IS

  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XINPUT
	PORT MAP (Z0 => Z0, XI0 => XI0);
END lattice_arch;
-- VHDL netlist for ID11
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ID11 IS 
    PORT (
        XI0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
END ID11;


ARCHITECTURE lattice_arch OF ID11 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI0);
END lattice_arch;
-- VHDL netlist for ID14
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ID14 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END ID14;


ARCHITECTURE lattice_arch OF ID14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : XINPUT
	PORT MAP (Z0 => UQVN_N2, XI0 => XI2);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, CLK => CLK);
UQVB_B6 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI1);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, CLK => CLK);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N4, XI0 => XI0);
END lattice_arch;
-- VHDL netlist for ID18
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ID18 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        XI4 : IN std_logic;
        XI5 : IN std_logic;
        XI6 : IN std_logic;
        XI7 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END ID18;


ARCHITECTURE lattice_arch OF ID18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, CLK => CLK);
UQVB_B4 : XINPUT
	PORT MAP (Z0 => UQVN_N2, XI0 => XI2);
UQVB_B5 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, CLK => CLK);
UQVB_B6 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI1);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, CLK => CLK);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N4, XI0 => XI0);
UQVB_B9 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N5, CLK => CLK);
UQVB_B10 : XINPUT
	PORT MAP (Z0 => UQVN_N5, XI0 => XI4);
UQVB_B11 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N6, CLK => CLK);
UQVB_B12 : XINPUT
	PORT MAP (Z0 => UQVN_N6, XI0 => XI5);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N7, CLK => CLK);
UQVB_B14 : XINPUT
	PORT MAP (Z0 => UQVN_N7, XI0 => XI6);
UQVB_B15 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N8, CLK => CLK);
UQVB_B16 : XINPUT
	PORT MAP (Z0 => UQVN_N8, XI0 => XI7);
END lattice_arch;
-- VHDL netlist for ID21
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ID21 IS 
    PORT (
        XI0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
END ID21;


ARCHITECTURE lattice_arch OF ID21 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, CLK => UQVN_N2);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
END lattice_arch;
-- VHDL netlist for ID24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ID24 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END ID24;


ARCHITECTURE lattice_arch OF ID24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => UQVN_N2);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N3, CLK => UQVN_N4);
UQVB_B5 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI2);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => CLK);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N5, CLK => UQVN_N6);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N5, XI0 => XI1);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => CLK);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N7, CLK => UQVN_N8);
UQVB_B11 : XINPUT
	PORT MAP (Z0 => UQVN_N7, XI0 => XI0);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => CLK);
END lattice_arch;
-- VHDL netlist for ID28
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY ID28 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        XI4 : IN std_logic;
        XI5 : IN std_logic;
        XI6 : IN std_logic;
        XI7 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END ID28;


ARCHITECTURE lattice_arch OF ID28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDFF1
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDFF1 use  entity  lat_vhd.XDFF1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XDFF1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, CLK => UQVN_N2);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => CLK);
UQVB_B4 : XDFF1
	PORT MAP (Q0 => Q2, D0 => UQVN_N3, CLK => UQVN_N4);
UQVB_B5 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI2);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => CLK);
UQVB_B7 : XDFF1
	PORT MAP (Q0 => Q1, D0 => UQVN_N5, CLK => UQVN_N6);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N5, XI0 => XI1);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => CLK);
UQVB_B10 : XDFF1
	PORT MAP (Q0 => Q0, D0 => UQVN_N7, CLK => UQVN_N8);
UQVB_B11 : XINPUT
	PORT MAP (Z0 => UQVN_N7, XI0 => XI0);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => CLK);
UQVB_B13 : XDFF1
	PORT MAP (Q0 => Q4, D0 => UQVN_N9, CLK => UQVN_N10);
UQVB_B14 : XINPUT
	PORT MAP (Z0 => UQVN_N9, XI0 => XI4);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => CLK);
UQVB_B16 : XDFF1
	PORT MAP (Q0 => Q5, D0 => UQVN_N11, CLK => UQVN_N12);
UQVB_B17 : XINPUT
	PORT MAP (Z0 => UQVN_N11, XI0 => XI5);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => CLK);
UQVB_B19 : XDFF1
	PORT MAP (Q0 => Q6, D0 => UQVN_N13, CLK => UQVN_N14);
UQVB_B20 : XINPUT
	PORT MAP (Z0 => UQVN_N13, XI0 => XI6);
UQVB_B21 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => CLK);
UQVB_B22 : XDFF1
	PORT MAP (Q0 => Q7, D0 => UQVN_N15, CLK => UQVN_N16);
UQVB_B23 : XINPUT
	PORT MAP (Z0 => UQVN_N15, XI0 => XI7);
UQVB_B24 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => CLK);
END lattice_arch;
-- VHDL netlist for IL11
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IL11 IS 
    PORT (
        XI0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
END IL11;


ARCHITECTURE lattice_arch OF IL11 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, G => G);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI0);
END lattice_arch;
-- VHDL netlist for IL14
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IL14 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END IL14;


ARCHITECTURE lattice_arch OF IL14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, G => G);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, G => G);
UQVB_B4 : XINPUT
	PORT MAP (Z0 => UQVN_N2, XI0 => XI2);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, G => G);
UQVB_B6 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI1);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, G => G);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N4, XI0 => XI0);
END lattice_arch;
-- VHDL netlist for IL18
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IL18 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        XI4 : IN std_logic;
        XI5 : IN std_logic;
        XI6 : IN std_logic;
        XI7 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END IL18;


ARCHITECTURE lattice_arch OF IL18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, G => G);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N2, G => G);
UQVB_B4 : XINPUT
	PORT MAP (Z0 => UQVN_N2, XI0 => XI2);
UQVB_B5 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N3, G => G);
UQVB_B6 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI1);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N4, G => G);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N4, XI0 => XI0);
UQVB_B9 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N5, G => G);
UQVB_B10 : XINPUT
	PORT MAP (Z0 => UQVN_N5, XI0 => XI4);
UQVB_B11 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N6, G => G);
UQVB_B12 : XINPUT
	PORT MAP (Z0 => UQVN_N6, XI0 => XI5);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N7, G => G);
UQVB_B14 : XINPUT
	PORT MAP (Z0 => UQVN_N7, XI0 => XI6);
UQVB_B15 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N8, G => G);
UQVB_B16 : XINPUT
	PORT MAP (Z0 => UQVN_N8, XI0 => XI7);
END lattice_arch;
-- VHDL netlist for IL21
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IL21 IS 
    PORT (
        XI0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
END IL21;


ARCHITECTURE lattice_arch OF IL21 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N1, G => UQVN_N2);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI0);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
END lattice_arch;
-- VHDL netlist for IL24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IL24 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END IL24;


ARCHITECTURE lattice_arch OF IL24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, G => UQVN_N2);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N3, G => UQVN_N4);
UQVB_B5 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI2);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N5, G => UQVN_N6);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N5, XI0 => XI1);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N7, G => UQVN_N8);
UQVB_B11 : XINPUT
	PORT MAP (Z0 => UQVN_N7, XI0 => XI0);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => G);
END lattice_arch;
-- VHDL netlist for IL28
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY IL28 IS 
    PORT (
        XI0 : IN std_logic;
        XI1 : IN std_logic;
        XI2 : IN std_logic;
        XI3 : IN std_logic;
        XI4 : IN std_logic;
        XI5 : IN std_logic;
        XI6 : IN std_logic;
        XI7 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END IL28;


ARCHITECTURE lattice_arch OF IL28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XDL1
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: XDL1 use  entity  lat_vhd.XDL1(lattice_arch);


  COMPONENT XINPUT
    PORT (
        XI0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XINPUT use  entity  lat_vhd.XINPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XDL1
	PORT MAP (Q0 => Q3, D0 => UQVN_N1, G => UQVN_N2);
UQVB_B2 : XINPUT
	PORT MAP (Z0 => UQVN_N1, XI0 => XI3);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => G);
UQVB_B4 : XDL1
	PORT MAP (Q0 => Q2, D0 => UQVN_N3, G => UQVN_N4);
UQVB_B5 : XINPUT
	PORT MAP (Z0 => UQVN_N3, XI0 => XI2);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B7 : XDL1
	PORT MAP (Q0 => Q1, D0 => UQVN_N5, G => UQVN_N6);
UQVB_B8 : XINPUT
	PORT MAP (Z0 => UQVN_N5, XI0 => XI1);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B10 : XDL1
	PORT MAP (Q0 => Q0, D0 => UQVN_N7, G => UQVN_N8);
UQVB_B11 : XINPUT
	PORT MAP (Z0 => UQVN_N7, XI0 => XI0);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => G);
UQVB_B13 : XDL1
	PORT MAP (Q0 => Q4, D0 => UQVN_N9, G => UQVN_N10);
UQVB_B14 : XINPUT
	PORT MAP (Z0 => UQVN_N9, XI0 => XI4);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => G);
UQVB_B16 : XDL1
	PORT MAP (Q0 => Q5, D0 => UQVN_N11, G => UQVN_N12);
UQVB_B17 : XINPUT
	PORT MAP (Z0 => UQVN_N11, XI0 => XI5);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => G);
UQVB_B19 : XDL1
	PORT MAP (Q0 => Q6, D0 => UQVN_N13, G => UQVN_N14);
UQVB_B20 : XINPUT
	PORT MAP (Z0 => UQVN_N13, XI0 => XI6);
UQVB_B21 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B22 : XDL1
	PORT MAP (Q0 => Q7, D0 => UQVN_N15, G => UQVN_N16);
UQVB_B23 : XINPUT
	PORT MAP (Z0 => UQVN_N15, XI0 => XI7);
UQVB_B24 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => G);
END lattice_arch;
-- VHDL netlist for LD11
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD11 IS 
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic
    );
END LD11;


ARCHITECTURE lattice_arch OF LD11 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, NUIB_S0, NUIB_S1 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B2 : SHFE
	PORT MAP (REF => G, DATA => D0);
NUIB_C1 : BUF
	PORT MAP (Z0 => NUIB_S0, A0 => D0);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => NUIB_S0);
NUIB_C2 : BUF
	PORT MAP (Z0 => NUIB_S1, A0 => G);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => NUIB_S0, A1 => NUIB_S1);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B7 : PW
	PORT MAP (PULSE => G);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
END lattice_arch;
-- VHDL netlist for LD14
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD14 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD14;


ARCHITECTURE lattice_arch OF LD14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B2 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B3A : BUF
	PORT MAP (Z0 => UQVN_N21, A0 => D3);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => UQVN_N21);
UQVB_B4A : BUF
	PORT MAP (Z0 => UQVN_N22, A0 => G);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N21, A1 => UQVN_N22);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B7 : PW
	PORT MAP (PULSE => G);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N5);
UQVB_B9 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N8);
UQVB_B10 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B11A : BUF
	PORT MAP (Z0 => UQVN_N23, A0 => D2);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N23);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N23, A1 => UQVN_N22);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N9);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => G);
UQVB_B15 : PW
	PORT MAP (PULSE => G);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N10);
UQVB_B17 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N12, A1 => UQVN_N11, A2 => UQVN_N13);
UQVB_B18 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B19A : BUF
	PORT MAP (Z0 => UQVN_N24, A0 => D1);
UQVB_B19 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N15, A1 => UQVN_N24);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N24, A1 => UQVN_N22);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N15, A1 => UQVN_N14);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B23 : PW
	PORT MAP (PULSE => G);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N15);
UQVB_B25 : OR3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N18);
UQVB_B26 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B27A : BUF
	PORT MAP (Z0 => UQVN_N25, A0 => D0);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N20, A1 => UQVN_N25);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N25, A1 => UQVN_N22);
UQVB_B29 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => G);
UQVB_B31 : PW
	PORT MAP (PULSE => G);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N20);
END lattice_arch;
-- VHDL netlist for LD18
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD18 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        G : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD18;


ARCHITECTURE lattice_arch OF LD18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B2 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B3A : BUF
	PORT MAP (Z0 => UQVN_N41, A0 => D3);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => UQVN_N41);
UQVB_B4A : BUF
	PORT MAP (Z0 => UQVN_N49, A0 => G);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N41, A1 => UQVN_N49);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B7 : PW
	PORT MAP (PULSE => G);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N5);
UQVB_B9 : OR3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N8);
UQVB_B10 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B11A : BUF
	PORT MAP (Z0 => UQVN_N42, A0 => D2);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N42);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N42, A1 => UQVN_N49);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N9);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => G);
UQVB_B15 : PW
	PORT MAP (PULSE => G);
UQVB_B16 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N10);
UQVB_B17 : OR3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N12, A1 => UQVN_N11, A2 => UQVN_N13);
UQVB_B18 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B19A : BUF
	PORT MAP (Z0 => UQVN_N43, A0 => D1);
UQVB_B19 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N15, A1 => UQVN_N43);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N43, A1 => UQVN_N49);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N15, A1 => UQVN_N14);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B23 : PW
	PORT MAP (PULSE => G);
UQVB_B24 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N15);
UQVB_B25 : OR3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N18);
UQVB_B26 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B27A : BUF
	PORT MAP (Z0 => UQVN_N44, A0 => D0);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N20, A1 => UQVN_N44);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N44, A1 => UQVN_N49);
UQVB_B29 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => G);
UQVB_B31 : PW
	PORT MAP (PULSE => G);
UQVB_B32 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N20);
UQVB_B33 : OR3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N22, A1 => UQVN_N21, A2 => UQVN_N23);
UQVB_B34 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B35A : BUF
	PORT MAP (Z0 => UQVN_N45, A0 => D4);
UQVB_B35 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N25, A1 => UQVN_N45);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N45, A1 => UQVN_N49);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N25, A1 => UQVN_N24);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => G);
UQVB_B39 : PW
	PORT MAP (PULSE => G);
UQVB_B40 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N25);
UQVB_B41 : OR3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N28);
UQVB_B42 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B43A : BUF
	PORT MAP (Z0 => UQVN_N46, A0 => D5);
UQVB_B43 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N30, A1 => UQVN_N46);
UQVB_B44 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N46, A1 => UQVN_N49);
UQVB_B45 : AND2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N30, A1 => UQVN_N29);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => G);
UQVB_B47 : PW
	PORT MAP (PULSE => G);
UQVB_B48 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N30);
UQVB_B49 : OR3
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N33);
UQVB_B50 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B51A : BUF
	PORT MAP (Z0 => UQVN_N47, A0 => D6);
UQVB_B51 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N35, A1 => UQVN_N47);
UQVB_B52 : AND2
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N47, A1 => UQVN_N49);
UQVB_B53 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N35, A1 => UQVN_N34);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => G);
UQVB_B55 : PW
	PORT MAP (PULSE => G);
UQVB_B56 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N35);
UQVB_B57 : OR3
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N38);
UQVB_B58 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B59A : BUF
	PORT MAP (Z0 => UQVN_N48, A0 => D7);
UQVB_B59 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N40, A1 => UQVN_N48);
UQVB_B60 : AND2
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N48, A1 => UQVN_N49);
UQVB_B61 : AND2
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N40, A1 => UQVN_N39);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => G);
UQVB_B63 : PW
	PORT MAP (PULSE => G);
UQVB_B64 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N40);
END lattice_arch;
-- VHDL netlist for LD21
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD21 IS 
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END LD21;


ARCHITECTURE lattice_arch OF LD21 IS
SIGNAL   UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
		 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B2A : BUF
	PORT MAP (Z0 => UQVN_N7, A0 => D0);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N7);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N5);
UQVB_B4A : BUF
	PORT MAP (Z0 => UQVN_N8, A0 => G);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N7, A1 => UQVN_N4, A2 => UQVN_N8);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B7 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B8 : PW
	PORT MAP (PULSE => G);
UQVB_B9 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B10 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N6);
END lattice_arch;
-- VHDL netlist for LD24
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD24 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        G : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD24;


ARCHITECTURE lattice_arch OF LD24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B2A : BUF	
	PORT MAP (Z0 => UQVN_N25, A0 => D3);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N25);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N5);
UQVB_B4A : BUF	
	PORT MAP (Z0 => UQVN_N29, A0 => G);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N25, A1 => UQVN_N4, A2 => UQVN_N29);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B7 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B8 : PW
	PORT MAP (PULSE => G);
UQVB_B9 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B10 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N6);
UQVB_B12 : OR3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9);
UQVB_B13A : BUF	
	PORT MAP (Z0 => UQVN_N26, A0 => D2);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N12, A1 => UQVN_N10, A2 => UQVN_N26);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N12, A1 => UQVN_N10, A2 => UQVN_N11);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N26, A1 => UQVN_N10, A2 => UQVN_N29);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CD);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B18 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B19 : PW
	PORT MAP (PULSE => G);
UQVB_B20 : SHFE
	PORT MAP (REF => UQVN_N10, DATA => G);
UQVB_B21 : PW
	PORT MAP (PULSE => UQVN_N10);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N12);
UQVB_B23 : OR3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N15);
UQVB_B24A : BUF	
	PORT MAP (Z0 => UQVN_N27, A0 => D1);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N18, A1 => UQVN_N16, A2 => UQVN_N27);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N18, A1 => UQVN_N16, A2 => UQVN_N17);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N27, A1 => UQVN_N16, A2 => UQVN_N29);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => CD);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => G);
UQVB_B29 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B30 : PW
	PORT MAP (PULSE => G);
UQVB_B31 : SHFE
	PORT MAP (REF => UQVN_N16, DATA => G);
UQVB_B32 : PW
	PORT MAP (PULSE => UQVN_N16);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N18);
UQVB_B34 : OR3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N21);
UQVB_B35A : BUF	
	PORT MAP (Z0 => UQVN_N28, A0 => D0);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N24, A1 => UQVN_N22, A2 => UQVN_N28);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N24, A1 => UQVN_N22, A2 => UQVN_N23);
UQVB_B37 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N28, A1 => UQVN_N22, A2 => UQVN_N29);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B40 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B41 : PW
	PORT MAP (PULSE => G);
UQVB_B42 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B43 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B44 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N24);
END lattice_arch;
-- VHDL netlist for LD28
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD28 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        G : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD28;


ARCHITECTURE lattice_arch OF LD28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B2A : BUF
	PORT MAP (Z0 => UQVN_N49, A0 => D3);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N49);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N5);
UQVB_B4A : BUF
	PORT MAP (Z0 => UQVN_N57, A0 => G);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N49, A1 => UQVN_N4, A2 => UQVN_N57);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B7 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B8 : PW
	PORT MAP (PULSE => G);
UQVB_B9 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B10 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N6);
UQVB_B12 : OR3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9);
UQVB_B13A : BUF
	PORT MAP (Z0 => UQVN_N50, A0 => D2);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N12, A1 => UQVN_N10, A2 => UQVN_N50);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N12, A1 => UQVN_N10, A2 => UQVN_N11);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N50, A1 => UQVN_N10, A2 => UQVN_N57);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CD);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B18 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B19 : PW
	PORT MAP (PULSE => G);
UQVB_B20 : SHFE
	PORT MAP (REF => UQVN_N10, DATA => G);
UQVB_B21 : PW
	PORT MAP (PULSE => UQVN_N10);
UQVB_B22 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N12);
UQVB_B23 : OR3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N15);
UQVB_B24A : BUF
	PORT MAP (Z0 => UQVN_N51, A0 => D1);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N18, A1 => UQVN_N16, A2 => UQVN_N51);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N18, A1 => UQVN_N16, A2 => UQVN_N17);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N51, A1 => UQVN_N16, A2 => UQVN_N57);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => CD);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => G);
UQVB_B29 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B30 : PW
	PORT MAP (PULSE => G);
UQVB_B31 : SHFE
	PORT MAP (REF => UQVN_N16, DATA => G);
UQVB_B32 : PW
	PORT MAP (PULSE => UQVN_N16);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N18);
UQVB_B34 : OR3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N21);
UQVB_B35A : BUF
	PORT MAP (Z0 => UQVN_N52, A0 => D0);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N24, A1 => UQVN_N22, A2 => UQVN_N52);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N24, A1 => UQVN_N22, A2 => UQVN_N23);
UQVB_B37 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N52, A1 => UQVN_N22, A2 => UQVN_N57);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B40 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B41 : PW
	PORT MAP (PULSE => G);
UQVB_B42 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B43 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B44 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N24);
UQVB_B45 : OR3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N27);
UQVB_B46A : BUF
	PORT MAP (Z0 => UQVN_N53, A0 => D6);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N30, A1 => UQVN_N28, A2 => UQVN_N53);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N30, A1 => UQVN_N28, A2 => UQVN_N29);
UQVB_B48 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N53, A1 => UQVN_N28, A2 => UQVN_N57);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => CD);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => G);
UQVB_B51 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B52 : PW
	PORT MAP (PULSE => G);
UQVB_B53 : SHFE
	PORT MAP (REF => UQVN_N28, DATA => G);
UQVB_B54 : PW
	PORT MAP (PULSE => UQVN_N28);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N30);
UQVB_B56 : OR3
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N33);
UQVB_B57A : BUF
	PORT MAP (Z0 => UQVN_N54, A0 => D5);
UQVB_B57 : AND3
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => UQVN_N34, A2 => UQVN_N54);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N36, A1 => UQVN_N34, A2 => UQVN_N35);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N54, A1 => UQVN_N34, A2 => UQVN_N57);
UQVB_B60 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => CD);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => G);
UQVB_B62 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B63 : PW
	PORT MAP (PULSE => G);
UQVB_B64 : SHFE
	PORT MAP (REF => UQVN_N34, DATA => G);
UQVB_B65 : PW
	PORT MAP (PULSE => UQVN_N34);
UQVB_B66 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N36);
UQVB_B67 : OR3
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N39);
UQVB_B68A : BUF
	PORT MAP (Z0 => UQVN_N55, A0 => D4);
UQVB_B68 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N42, A1 => UQVN_N40, A2 => UQVN_N55);
UQVB_B69 : AND3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N42, A1 => UQVN_N40, A2 => UQVN_N41);
UQVB_B70 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N55, A1 => UQVN_N40, A2 => UQVN_N57);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CD);
UQVB_B72 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => G);
UQVB_B73 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B74 : PW
	PORT MAP (PULSE => G);
UQVB_B75 : SHFE
	PORT MAP (REF => UQVN_N40, DATA => G);
UQVB_B76 : PW
	PORT MAP (PULSE => UQVN_N40);
UQVB_B77 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N42);
UQVB_B78 : OR3
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N44, A1 => UQVN_N43, A2 => UQVN_N45);
UQVB_B79A : BUF
	PORT MAP (Z0 => UQVN_N56, A0 => D7);
UQVB_B79 : AND3
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N48, A1 => UQVN_N46, A2 => UQVN_N56);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N48, A1 => UQVN_N46, A2 => UQVN_N47);
UQVB_B81 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N56, A1 => UQVN_N46, A2 => UQVN_N57);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => CD);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => G);
UQVB_B84 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B85 : PW
	PORT MAP (PULSE => G);
UQVB_B86 : SHFE
	PORT MAP (REF => UQVN_N46, DATA => G);
UQVB_B87 : PW
	PORT MAP (PULSE => UQVN_N46);
UQVB_B88 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N48);
END lattice_arch;
-- VHDL netlist for LD31
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD31 IS 
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        Q0 : OUT std_logic
    );
END LD31;


ARCHITECTURE lattice_arch OF LD31 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
		 UQVN_N5, UQVN_N6, UQVN_N7 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => PD);
UQVB_B2A0 : BUF
	PORT MAP (Z0 => UQVN_N6, A0 => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B4A0 : BUF
	PORT MAP (Z0 => UQVN_N7, A0 => G);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N6, A1 => UQVN_N7);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B6 : PW
	PORT MAP (PULSE => G);
UQVB_B7 : PW
	PORT MAP (PULSE => PD);
UQVB_B8 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B9 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
END lattice_arch;
-- VHDL netlist for LD34
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD34;


ARCHITECTURE lattice_arch OF LD34 IS
SIGNAL UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
 	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => PD);
UQVB_B2A : BUF
	PORT MAP (Z0 => UQVN_N21, A0 => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => UQVN_N21);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B4A : BUF
	PORT MAP (Z0 => UQVN_N25, A0 => G);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N21, A1 => UQVN_N25);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B6 : PW
	PORT MAP (PULSE => G);
UQVB_B7 : PW
	PORT MAP (PULSE => PD);
UQVB_B8 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B9 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N5);
UQVB_B11 : OR4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N8, 
	A3 => PD);
UQVB_B12A : BUF
	PORT MAP (Z0 => UQVN_N23, A0 => D2);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N23);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N9);
UQVB_B14 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N23, A1 => UQVN_N25);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => G);
UQVB_B16 : PW
	PORT MAP (PULSE => G);
UQVB_B17 : PW
	PORT MAP (PULSE => PD);
UQVB_B18 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B19 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N10);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N12, A1 => UQVN_N11, A2 => UQVN_N13, 
	A3 => PD);
UQVB_B22A : BUF
	PORT MAP (Z0 => UQVN_N24, A0 => D1);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N15, A1 => UQVN_N24);
UQVB_B23 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N15, A1 => UQVN_N14);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N24, A1 => UQVN_N25);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B26 : PW
	PORT MAP (PULSE => G);
UQVB_B27 : PW
	PORT MAP (PULSE => PD);
UQVB_B28 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B29 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N15);
UQVB_B31 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N18, 
	A3 => PD);
UQVB_B32A : BUF
	PORT MAP (Z0 => UQVN_N22, A0 => D0);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N20, A1 => UQVN_N22);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N22, A1 => UQVN_N25);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => G);
UQVB_B36 : PW
	PORT MAP (PULSE => G);
UQVB_B37 : PW
	PORT MAP (PULSE => PD);
UQVB_B38 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B39 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B40 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N20);
END lattice_arch;
-- VHDL netlist for LD38
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD38;


ARCHITECTURE lattice_arch OF LD38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => PD);
UQVB_B2A : BUF
	PORT MAP (Z0 => UQVN_N41, A0 => D7);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => UQVN_N41);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B4A : BUF
	PORT MAP (Z0 => UQVN_N49, A0 => G);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N41, A1 => UQVN_N49);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B6 : PW
	PORT MAP (PULSE => G);
UQVB_B7 : PW
	PORT MAP (PULSE => PD);
UQVB_B8 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B9 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N5);
UQVB_B11 : OR4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N8, 
	A3 => PD);
UQVB_B11A : BUF
	PORT MAP (Z0 => UQVN_N42, A0 => D6);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N42);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N9);
UQVB_B14 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N42, A1 => UQVN_N49);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => G);
UQVB_B16 : PW
	PORT MAP (PULSE => G);
UQVB_B17 : PW
	PORT MAP (PULSE => PD);
UQVB_B18 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B19 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B20 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N10);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N12, A1 => UQVN_N11, A2 => UQVN_N13, 
	A3 => PD);
UQVB_B19A : BUF
	PORT MAP (Z0 => UQVN_N43, A0 => D5);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N15, A1 => UQVN_N43);
UQVB_B23 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N15, A1 => UQVN_N14);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N43, A1 => UQVN_N49);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B26 : PW
	PORT MAP (PULSE => G);
UQVB_B27 : PW
	PORT MAP (PULSE => PD);
UQVB_B28 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B29 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N15);
UQVB_B31 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N18, 
	A3 => PD);
UQVB_B35A : BUF
	PORT MAP (Z0 => UQVN_N45, A0 => D4);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N20, A1 => UQVN_N45);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N45, A1 => UQVN_N49);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => G);
UQVB_B36 : PW
	PORT MAP (PULSE => G);
UQVB_B37 : PW
	PORT MAP (PULSE => PD);
UQVB_B38 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B39 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B40 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N20);
UQVB_B41 : OR4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N22, A1 => UQVN_N21, A2 => UQVN_N23, 
	A3 => PD);
UQVB_B27A : BUF
	PORT MAP (Z0 => UQVN_N44, A0 => D2);
UQVB_B42 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N25, A1 => UQVN_N44);
UQVB_B43 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N25, A1 => UQVN_N24);
UQVB_B44 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N44, A1 => UQVN_N44);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => G);
UQVB_B46 : PW
	PORT MAP (PULSE => G);
UQVB_B47 : PW
	PORT MAP (PULSE => PD);
UQVB_B48 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B49 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B50 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N25);
UQVB_B51 : OR4
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N28, 
	A3 => PD);
UQVB_B43A : BUF
	PORT MAP (Z0 => UQVN_N46, A0 => D3);
UQVB_B52 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N30, A1 => UQVN_N46);
UQVB_B53 : AND2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N30, A1 => UQVN_N29);
UQVB_B54 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N46, A1 => UQVN_N46);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => G);
UQVB_B56 : PW
	PORT MAP (PULSE => G);
UQVB_B57 : PW
	PORT MAP (PULSE => PD);
UQVB_B58 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B59 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B60 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N30);
UQVB_B61 : OR4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N33, 
	A3 => PD);
UQVB_B51A : BUF
	PORT MAP (Z0 => UQVN_N47, A0 => D1);
UQVB_B62 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N35, A1 => UQVN_N47);
UQVB_B63 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N35, A1 => UQVN_N34);
UQVB_B64 : AND2
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N47, A1 => UQVN_N49);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => G);
UQVB_B66 : PW
	PORT MAP (PULSE => G);
UQVB_B67 : PW
	PORT MAP (PULSE => PD);
UQVB_B68 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B69 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B70 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N35);
UQVB_B71 : OR4
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N38, 
	A3 => PD);
UQVB_B59A : BUF
	PORT MAP (Z0 => UQVN_N48, A0 => D0);
UQVB_B72 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N40, A1 => UQVN_N48);
UQVB_B73 : AND2
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N40, A1 => UQVN_N39);
UQVB_B74 : AND2
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N48, A1 => UQVN_N49);
UQVB_B75 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => G);
UQVB_B76 : PW
	PORT MAP (PULSE => G);
UQVB_B77 : PW
	PORT MAP (PULSE => PD);
UQVB_B78 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B79 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B80 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N40);
END lattice_arch;
-- VHDL netlist for LD41
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD41 IS 
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END LD41;


ARCHITECTURE lattice_arch OF LD41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N7, A1 => UQVN_N4, A2 => D0);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N7, A1 => UQVN_N4, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => UQVN_N4, A2 => G);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N4, A1 => PD);
UQVB_B6 : OR4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => UQVN_N5);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B8 : PW
	PORT MAP (PULSE => G);
UQVB_B9 : PW
	PORT MAP (PULSE => PD);
UQVB_B10 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B11 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B12 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B13 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N7);
UQVB_B15 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => PD);
END lattice_arch;
-- VHDL netlist for LD44
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD44;


ARCHITECTURE lattice_arch OF LD44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N7, A1 => UQVN_N4, A2 => D3);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N7, A1 => UQVN_N4, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => UQVN_N4, A2 => G);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N4, A1 => PD);
UQVB_B6 : OR4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => UQVN_N5);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B8 : PW
	PORT MAP (PULSE => G);
UQVB_B9 : PW
	PORT MAP (PULSE => PD);
UQVB_B10 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B11 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B12 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B13 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N7);
UQVB_B15 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => PD);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => CD);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N14, A1 => UQVN_N11, A2 => D2);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N14, A1 => UQVN_N11, A2 => UQVN_N13);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D2, A1 => UQVN_N11, A2 => G);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N11, A1 => PD);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N9, A1 => UQVN_N8, A2 => UQVN_N10, 
	A3 => UQVN_N12);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => G);
UQVB_B23 : PW
	PORT MAP (PULSE => G);
UQVB_B24 : PW
	PORT MAP (PULSE => PD);
UQVB_B25 : PW
	PORT MAP (PULSE => UQVN_N11);
UQVB_B26 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => G);
UQVB_B27 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B28 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N14);
UQVB_B30 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => PD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => CD);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N21, A1 => UQVN_N18, A2 => D1);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => UQVN_N18, A2 => UQVN_N20);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => D1, A1 => UQVN_N18, A2 => G);
UQVB_B35 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N18, A1 => PD);
UQVB_B36 : OR4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N16, A1 => UQVN_N15, A2 => UQVN_N17, 
	A3 => UQVN_N19);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => G);
UQVB_B38 : PW
	PORT MAP (PULSE => G);
UQVB_B39 : PW
	PORT MAP (PULSE => PD);
UQVB_B40 : PW
	PORT MAP (PULSE => UQVN_N18);
UQVB_B41 : SHFE
	PORT MAP (REF => UQVN_N18, DATA => G);
UQVB_B42 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B43 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B44 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N21);
UQVB_B45 : SHFE
	PORT MAP (REF => UQVN_N18, DATA => PD);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => CD);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N28, A1 => UQVN_N25, A2 => D0);
UQVB_B48 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N28, A1 => UQVN_N25, A2 => UQVN_N27);
UQVB_B49 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => D0, A1 => UQVN_N25, A2 => G);
UQVB_B50 : AND2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N25, A1 => PD);
UQVB_B51 : OR4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N23, A1 => UQVN_N22, A2 => UQVN_N24, 
	A3 => UQVN_N26);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => G);
UQVB_B53 : PW
	PORT MAP (PULSE => G);
UQVB_B54 : PW
	PORT MAP (PULSE => PD);
UQVB_B55 : PW
	PORT MAP (PULSE => UQVN_N25);
UQVB_B56 : SHFE
	PORT MAP (REF => UQVN_N25, DATA => G);
UQVB_B57 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B58 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B59 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N28);
UQVB_B60 : SHFE
	PORT MAP (REF => UQVN_N25, DATA => PD);
END lattice_arch;
-- VHDL netlist for LD48
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD48;


ARCHITECTURE lattice_arch OF LD48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N7, A1 => UQVN_N4, A2 => D3);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N7, A1 => UQVN_N4, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => UQVN_N4, A2 => G);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N4, A1 => PD);
UQVB_B6 : OR4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => UQVN_N5);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => G);
UQVB_B8 : PW
	PORT MAP (PULSE => G);
UQVB_B9 : PW
	PORT MAP (PULSE => PD);
UQVB_B10 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B11 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B12 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B13 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B14 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N7);
UQVB_B15 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => PD);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => CD);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N14, A1 => UQVN_N11, A2 => D2);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N14, A1 => UQVN_N11, A2 => UQVN_N13);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D2, A1 => UQVN_N11, A2 => G);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N11, A1 => PD);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N9, A1 => UQVN_N8, A2 => UQVN_N10, 
	A3 => UQVN_N12);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => G);
UQVB_B23 : PW
	PORT MAP (PULSE => G);
UQVB_B24 : PW
	PORT MAP (PULSE => PD);
UQVB_B25 : PW
	PORT MAP (PULSE => UQVN_N11);
UQVB_B26 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => G);
UQVB_B27 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B28 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N14);
UQVB_B30 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => PD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => CD);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N21, A1 => UQVN_N18, A2 => D1);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => UQVN_N18, A2 => UQVN_N20);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => D1, A1 => UQVN_N18, A2 => G);
UQVB_B35 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N18, A1 => PD);
UQVB_B36 : OR4
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N16, A1 => UQVN_N15, A2 => UQVN_N17, 
	A3 => UQVN_N19);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => G);
UQVB_B38 : PW
	PORT MAP (PULSE => G);
UQVB_B39 : PW
	PORT MAP (PULSE => PD);
UQVB_B40 : PW
	PORT MAP (PULSE => UQVN_N18);
UQVB_B41 : SHFE
	PORT MAP (REF => UQVN_N18, DATA => G);
UQVB_B42 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B43 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B44 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N21);
UQVB_B45 : SHFE
	PORT MAP (REF => UQVN_N18, DATA => PD);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => CD);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N28, A1 => UQVN_N25, A2 => D0);
UQVB_B48 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N28, A1 => UQVN_N25, A2 => UQVN_N27);
UQVB_B49 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => D0, A1 => UQVN_N25, A2 => G);
UQVB_B50 : AND2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N25, A1 => PD);
UQVB_B51 : OR4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N23, A1 => UQVN_N22, A2 => UQVN_N24, 
	A3 => UQVN_N26);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => G);
UQVB_B53 : PW
	PORT MAP (PULSE => G);
UQVB_B54 : PW
	PORT MAP (PULSE => PD);
UQVB_B55 : PW
	PORT MAP (PULSE => UQVN_N25);
UQVB_B56 : SHFE
	PORT MAP (REF => UQVN_N25, DATA => G);
UQVB_B57 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B58 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B59 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N28);
UQVB_B60 : SHFE
	PORT MAP (REF => UQVN_N25, DATA => PD);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => CD);
UQVB_B62 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N35, A1 => UQVN_N32, A2 => D7);
UQVB_B63 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N35, A1 => UQVN_N32, A2 => UQVN_N34);
UQVB_B64 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => D7, A1 => UQVN_N32, A2 => G);
UQVB_B65 : AND2
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N32, A1 => PD);
UQVB_B66 : OR4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N30, A1 => UQVN_N29, A2 => UQVN_N31, 
	A3 => UQVN_N33);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => G);
UQVB_B68 : PW
	PORT MAP (PULSE => G);
UQVB_B69 : PW
	PORT MAP (PULSE => PD);
UQVB_B70 : PW
	PORT MAP (PULSE => UQVN_N32);
UQVB_B71 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => G);
UQVB_B72 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B73 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B74 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N35);
UQVB_B75 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => PD);
UQVB_B76 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => CD);
UQVB_B77 : AND3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N42, A1 => UQVN_N39, A2 => D6);
UQVB_B78 : AND3
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N42, A1 => UQVN_N39, A2 => UQVN_N41);
UQVB_B79 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => D6, A1 => UQVN_N39, A2 => G);
UQVB_B80 : AND2
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N39, A1 => PD);
UQVB_B81 : OR4
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N38, 
	A3 => UQVN_N40);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => G);
UQVB_B83 : PW
	PORT MAP (PULSE => G);
UQVB_B84 : PW
	PORT MAP (PULSE => PD);
UQVB_B85 : PW
	PORT MAP (PULSE => UQVN_N39);
UQVB_B86 : SHFE
	PORT MAP (REF => UQVN_N39, DATA => G);
UQVB_B87 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B88 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B89 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N42);
UQVB_B90 : SHFE
	PORT MAP (REF => UQVN_N39, DATA => PD);
UQVB_B91 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => CD);
UQVB_B92 : AND3
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N49, A1 => UQVN_N46, A2 => D5);
UQVB_B93 : AND3
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N49, A1 => UQVN_N46, A2 => UQVN_N48);
UQVB_B94 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => D5, A1 => UQVN_N46, A2 => G);
UQVB_B95 : AND2
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N46, A1 => PD);
UQVB_B96 : OR4
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N44, A1 => UQVN_N43, A2 => UQVN_N45, 
	A3 => UQVN_N47);
UQVB_B97 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => G);
UQVB_B98 : PW
	PORT MAP (PULSE => G);
UQVB_B99 : PW
	PORT MAP (PULSE => PD);
UQVB_B100 : PW
	PORT MAP (PULSE => UQVN_N46);
UQVB_B101 : SHFE
	PORT MAP (REF => UQVN_N46, DATA => G);
UQVB_B102 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B103 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B104 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N49);
UQVB_B105 : SHFE
	PORT MAP (REF => UQVN_N46, DATA => PD);
UQVB_B106 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => CD);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N56, A1 => UQVN_N53, A2 => D4);
UQVB_B108 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N56, A1 => UQVN_N53, A2 => UQVN_N55);
UQVB_B109 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => D4, A1 => UQVN_N53, A2 => G);
UQVB_B110 : AND2
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N53, A1 => PD);
UQVB_B111 : OR4
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N51, A1 => UQVN_N50, A2 => UQVN_N52, 
	A3 => UQVN_N54);
UQVB_B112 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => G);
UQVB_B113 : PW
	PORT MAP (PULSE => G);
UQVB_B114 : PW
	PORT MAP (PULSE => PD);
UQVB_B115 : PW
	PORT MAP (PULSE => UQVN_N53);
UQVB_B116 : SHFE
	PORT MAP (REF => UQVN_N53, DATA => G);
UQVB_B117 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B118 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B119 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N56);
UQVB_B120 : SHFE
	PORT MAP (REF => UQVN_N53, DATA => PD);
END lattice_arch;
-- VHDL netlist for LD51
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD51 IS 
    PORT (
        D0 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END LD51;


ARCHITECTURE lattice_arch OF LD51 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => PD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => D0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N5);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => UQVN_N4, A2 => G);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B8 : PW
	PORT MAP (PULSE => PD);
UQVB_B9 : PW
	PORT MAP (PULSE => G);
UQVB_B10 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B11 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B12 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N6);
UQVB_B14 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => PD);
END lattice_arch;
-- VHDL netlist for LD54
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD54 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD54;


ARCHITECTURE lattice_arch OF LD54 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => PD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => D3);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N5);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => UQVN_N4, A2 => G);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B8 : PW
	PORT MAP (PULSE => PD);
UQVB_B9 : PW
	PORT MAP (PULSE => G);
UQVB_B10 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B11 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B12 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N6);
UQVB_B14 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => PD);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CD);
UQVB_B16 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9, 
	A3 => PD);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N12, A1 => UQVN_N10, A2 => D2);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N12, A1 => UQVN_N10, A2 => UQVN_N11);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => D2, A1 => UQVN_N10, A2 => G);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B21 : PW
	PORT MAP (PULSE => UQVN_N10);
UQVB_B22 : PW
	PORT MAP (PULSE => PD);
UQVB_B23 : PW
	PORT MAP (PULSE => G);
UQVB_B24 : SHFE
	PORT MAP (REF => UQVN_N10, DATA => G);
UQVB_B25 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B26 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N12);
UQVB_B28 : SHFE
	PORT MAP (REF => UQVN_N10, DATA => PD);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => CD);
UQVB_B30 : OR4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N15, 
	A3 => PD);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N18, A1 => UQVN_N16, A2 => D1);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N18, A1 => UQVN_N16, A2 => UQVN_N17);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => D1, A1 => UQVN_N16, A2 => G);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => G);
UQVB_B35 : PW
	PORT MAP (PULSE => UQVN_N16);
UQVB_B36 : PW
	PORT MAP (PULSE => PD);
UQVB_B37 : PW
	PORT MAP (PULSE => G);
UQVB_B38 : SHFE
	PORT MAP (REF => UQVN_N16, DATA => G);
UQVB_B39 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B40 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B41 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N18);
UQVB_B42 : SHFE
	PORT MAP (REF => UQVN_N16, DATA => PD);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B44 : OR4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N21, 
	A3 => PD);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N24, A1 => UQVN_N22, A2 => D0);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N24, A1 => UQVN_N22, A2 => UQVN_N23);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D0, A1 => UQVN_N22, A2 => G);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B49 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B50 : PW
	PORT MAP (PULSE => PD);
UQVB_B51 : PW
	PORT MAP (PULSE => G);
UQVB_B52 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B53 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B54 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N24);
UQVB_B56 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => PD);
END lattice_arch;
-- VHDL netlist for LD58
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD58 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD58;


ARCHITECTURE lattice_arch OF LD58 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3, 
	A3 => PD);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => D3);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N5);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => UQVN_N4, A2 => G);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B8 : PW
	PORT MAP (PULSE => PD);
UQVB_B9 : PW
	PORT MAP (PULSE => G);
UQVB_B10 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B11 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B12 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B13 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N6);
UQVB_B14 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => PD);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CD);
UQVB_B16 : OR4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9, 
	A3 => PD);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N12, A1 => UQVN_N10, A2 => D2);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N12, A1 => UQVN_N10, A2 => UQVN_N11);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => D2, A1 => UQVN_N10, A2 => G);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => G);
UQVB_B21 : PW
	PORT MAP (PULSE => UQVN_N10);
UQVB_B22 : PW
	PORT MAP (PULSE => PD);
UQVB_B23 : PW
	PORT MAP (PULSE => G);
UQVB_B24 : SHFE
	PORT MAP (REF => UQVN_N10, DATA => G);
UQVB_B25 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B26 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N12);
UQVB_B28 : SHFE
	PORT MAP (REF => UQVN_N10, DATA => PD);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => CD);
UQVB_B30 : OR4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N15, 
	A3 => PD);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N18, A1 => UQVN_N16, A2 => D1);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N18, A1 => UQVN_N16, A2 => UQVN_N17);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => D1, A1 => UQVN_N16, A2 => G);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => G);
UQVB_B35 : PW
	PORT MAP (PULSE => UQVN_N16);
UQVB_B36 : PW
	PORT MAP (PULSE => PD);
UQVB_B37 : PW
	PORT MAP (PULSE => G);
UQVB_B38 : SHFE
	PORT MAP (REF => UQVN_N16, DATA => G);
UQVB_B39 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B40 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B41 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N18);
UQVB_B42 : SHFE
	PORT MAP (REF => UQVN_N16, DATA => PD);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B44 : OR4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N21, 
	A3 => PD);
UQVB_B45 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N24, A1 => UQVN_N22, A2 => D0);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N24, A1 => UQVN_N22, A2 => UQVN_N23);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D0, A1 => UQVN_N22, A2 => G);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B49 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B50 : PW
	PORT MAP (PULSE => PD);
UQVB_B51 : PW
	PORT MAP (PULSE => G);
UQVB_B52 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B53 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B54 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N24);
UQVB_B56 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => PD);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => CD);
UQVB_B58 : OR4
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N27, 
	A3 => PD);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N30, A1 => UQVN_N28, A2 => D7);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N30, A1 => UQVN_N28, A2 => UQVN_N29);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => D7, A1 => UQVN_N28, A2 => G);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => G);
UQVB_B63 : PW
	PORT MAP (PULSE => UQVN_N28);
UQVB_B64 : PW
	PORT MAP (PULSE => PD);
UQVB_B65 : PW
	PORT MAP (PULSE => G);
UQVB_B66 : SHFE
	PORT MAP (REF => UQVN_N28, DATA => G);
UQVB_B67 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B68 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B69 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N30);
UQVB_B70 : SHFE
	PORT MAP (REF => UQVN_N28, DATA => PD);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => CD);
UQVB_B72 : OR4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N33, 
	A3 => PD);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => UQVN_N34, A2 => D6);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N36, A1 => UQVN_N34, A2 => UQVN_N35);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => D6, A1 => UQVN_N34, A2 => G);
UQVB_B76 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => G);
UQVB_B77 : PW
	PORT MAP (PULSE => UQVN_N34);
UQVB_B78 : PW
	PORT MAP (PULSE => PD);
UQVB_B79 : PW
	PORT MAP (PULSE => G);
UQVB_B80 : SHFE
	PORT MAP (REF => UQVN_N34, DATA => G);
UQVB_B81 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B82 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B83 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N36);
UQVB_B84 : SHFE
	PORT MAP (REF => UQVN_N34, DATA => PD);
UQVB_B85 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CD);
UQVB_B86 : OR4
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N39, 
	A3 => PD);
UQVB_B87 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N42, A1 => UQVN_N40, A2 => D5);
UQVB_B88 : AND3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N42, A1 => UQVN_N40, A2 => UQVN_N41);
UQVB_B89 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => D5, A1 => UQVN_N40, A2 => G);
UQVB_B90 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => G);
UQVB_B91 : PW
	PORT MAP (PULSE => UQVN_N40);
UQVB_B92 : PW
	PORT MAP (PULSE => PD);
UQVB_B93 : PW
	PORT MAP (PULSE => G);
UQVB_B94 : SHFE
	PORT MAP (REF => UQVN_N40, DATA => G);
UQVB_B95 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B96 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B97 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N42);
UQVB_B98 : SHFE
	PORT MAP (REF => UQVN_N40, DATA => PD);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => CD);
UQVB_B100 : OR4
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N44, A1 => UQVN_N43, A2 => UQVN_N45, 
	A3 => PD);
UQVB_B101 : AND3
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N48, A1 => UQVN_N46, A2 => D4);
UQVB_B102 : AND3
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N48, A1 => UQVN_N46, A2 => UQVN_N47);
UQVB_B103 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => D4, A1 => UQVN_N46, A2 => G);
UQVB_B104 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => G);
UQVB_B105 : PW
	PORT MAP (PULSE => UQVN_N46);
UQVB_B106 : PW
	PORT MAP (PULSE => PD);
UQVB_B107 : PW
	PORT MAP (PULSE => G);
UQVB_B108 : SHFE
	PORT MAP (REF => UQVN_N46, DATA => G);
UQVB_B109 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B110 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B111 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N48);
UQVB_B112 : SHFE
	PORT MAP (REF => UQVN_N46, DATA => PD);
END lattice_arch;
-- VHDL netlist for LD61
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD61 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        G : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic
    );
END LD61;


ARCHITECTURE lattice_arch OF LD61 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => G);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B4 : PW
	PORT MAP (PULSE => G);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N8);
UQVB_B6 : OR5
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N2, A1 => UQVN_N5, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI0, A1 => TG);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N8, A1 => UQVN_N7, A2 => TI0);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N6, A2 => D0);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => TG);
UQVB_B12 : PW
	PORT MAP (PULSE => TG);
UQVB_B13 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
END lattice_arch;
-- VHDL netlist for LD64
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD64 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        G : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD64;


ARCHITECTURE lattice_arch OF LD64 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => G);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B4 : PW
	PORT MAP (PULSE => G);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N8);
UQVB_B6 : OR5
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N2, A1 => UQVN_N5, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TG);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N8, A1 => UQVN_N7, A2 => TI3);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N6, A2 => D3);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => TG);
UQVB_B12 : PW
	PORT MAP (PULSE => TG);
UQVB_B13 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B14 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => D2, A1 => G);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => G);
UQVB_B17 : PW
	PORT MAP (PULSE => G);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N16);
UQVB_B19 : OR5
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N10, A1 => UQVN_N13, A2 => UQVN_N9, 
	A3 => UQVN_N12, A4 => UQVN_N11);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI2, A1 => TG);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N16, A1 => UQVN_N15, A2 => UQVN_N14);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N16, A1 => UQVN_N15, A2 => TI2);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N16, A1 => UQVN_N14, A2 => D2);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => TG);
UQVB_B25 : PW
	PORT MAP (PULSE => TG);
UQVB_B26 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B27 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D1, A1 => G);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B30 : PW
	PORT MAP (PULSE => G);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N24);
UQVB_B32 : OR5
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N18, A1 => UQVN_N21, A2 => UQVN_N17, 
	A3 => UQVN_N20, A4 => UQVN_N19);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => TI1, A1 => TG);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N22);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N24, A1 => UQVN_N23, A2 => TI1);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N24, A1 => UQVN_N22, A2 => D1);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => TG);
UQVB_B38 : PW
	PORT MAP (PULSE => TG);
UQVB_B39 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B40 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B41 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => D0, A1 => G);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => G);
UQVB_B43 : PW
	PORT MAP (PULSE => G);
UQVB_B44 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N32);
UQVB_B45 : OR5
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N26, A1 => UQVN_N29, A2 => UQVN_N25, 
	A3 => UQVN_N28, A4 => UQVN_N27);
UQVB_B46 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => TI0, A1 => TG);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30);
UQVB_B48 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N32, A1 => UQVN_N31, A2 => TI0);
UQVB_B49 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N32, A1 => UQVN_N30, A2 => D0);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => TG);
UQVB_B51 : PW
	PORT MAP (PULSE => TG);
UQVB_B52 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
END lattice_arch;
-- VHDL netlist for LD68
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD68 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        G : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD68;


ARCHITECTURE lattice_arch OF LD68 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64 : std_logic;


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => G);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => G);
UQVB_B4 : PW
	PORT MAP (PULSE => G);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N8);
UQVB_B6 : OR5
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N2, A1 => UQVN_N5, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => TG);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N8, A1 => UQVN_N7, A2 => TI3);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N6, A2 => D3);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => TG);
UQVB_B12 : PW
	PORT MAP (PULSE => TG);
UQVB_B13 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B14 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => D2, A1 => G);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => G);
UQVB_B17 : PW
	PORT MAP (PULSE => G);
UQVB_B18 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N16);
UQVB_B19 : OR5
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N10, A1 => UQVN_N13, A2 => UQVN_N9, 
	A3 => UQVN_N12, A4 => UQVN_N11);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => TI2, A1 => TG);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N16, A1 => UQVN_N15, A2 => UQVN_N14);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N16, A1 => UQVN_N15, A2 => TI2);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N16, A1 => UQVN_N14, A2 => D2);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => TG);
UQVB_B25 : PW
	PORT MAP (PULSE => TG);
UQVB_B26 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B27 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D1, A1 => G);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B30 : PW
	PORT MAP (PULSE => G);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N24);
UQVB_B32 : OR5
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N18, A1 => UQVN_N21, A2 => UQVN_N17, 
	A3 => UQVN_N20, A4 => UQVN_N19);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => TI1, A1 => TG);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N22);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N24, A1 => UQVN_N23, A2 => TI1);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N24, A1 => UQVN_N22, A2 => D1);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => TG);
UQVB_B38 : PW
	PORT MAP (PULSE => TG);
UQVB_B39 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B40 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B41 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => D0, A1 => G);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => G);
UQVB_B43 : PW
	PORT MAP (PULSE => G);
UQVB_B44 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N32);
UQVB_B45 : OR5
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N26, A1 => UQVN_N29, A2 => UQVN_N25, 
	A3 => UQVN_N28, A4 => UQVN_N27);
UQVB_B46 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => TI0, A1 => TG);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N32, A1 => UQVN_N31, A2 => UQVN_N30);
UQVB_B48 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N32, A1 => UQVN_N31, A2 => TI0);
UQVB_B49 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N32, A1 => UQVN_N30, A2 => D0);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => TG);
UQVB_B51 : PW
	PORT MAP (PULSE => TG);
UQVB_B52 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B53 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B54 : AND2
	PORT MAP (Z0 => UQVN_N35, A0 => D6, A1 => G);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => G);
UQVB_B56 : PW
	PORT MAP (PULSE => G);
UQVB_B57 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N40);
UQVB_B58 : OR5
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N34, A1 => UQVN_N37, A2 => UQVN_N33, 
	A3 => UQVN_N36, A4 => UQVN_N35);
UQVB_B59 : AND2
	PORT MAP (Z0 => UQVN_N36, A0 => TI6, A1 => TG);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N39, A2 => UQVN_N38);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N40, A1 => UQVN_N39, A2 => TI6);
UQVB_B62 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N40, A1 => UQVN_N38, A2 => D6);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => TG);
UQVB_B64 : PW
	PORT MAP (PULSE => TG);
UQVB_B65 : SHFE
	PORT MAP (REF => TG, DATA => TI6);
UQVB_B66 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B67 : AND2
	PORT MAP (Z0 => UQVN_N43, A0 => D5, A1 => G);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => G);
UQVB_B69 : PW
	PORT MAP (PULSE => G);
UQVB_B70 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N48);
UQVB_B71 : OR5
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N42, A1 => UQVN_N45, A2 => UQVN_N41, 
	A3 => UQVN_N44, A4 => UQVN_N43);
UQVB_B72 : AND2
	PORT MAP (Z0 => UQVN_N44, A0 => TI5, A1 => TG);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N48, A1 => UQVN_N47, A2 => UQVN_N46);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N48, A1 => UQVN_N47, A2 => TI5);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N48, A1 => UQVN_N46, A2 => D5);
UQVB_B76 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => TG);
UQVB_B77 : PW
	PORT MAP (PULSE => TG);
UQVB_B78 : SHFE
	PORT MAP (REF => TG, DATA => TI5);
UQVB_B79 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B80 : AND2
	PORT MAP (Z0 => UQVN_N51, A0 => D4, A1 => G);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => G);
UQVB_B82 : PW
	PORT MAP (PULSE => G);
UQVB_B83 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N56);
UQVB_B84 : OR5
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N50, A1 => UQVN_N53, A2 => UQVN_N49, 
	A3 => UQVN_N52, A4 => UQVN_N51);
UQVB_B85 : AND2
	PORT MAP (Z0 => UQVN_N52, A0 => TI4, A1 => TG);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N56, A1 => UQVN_N55, A2 => UQVN_N54);
UQVB_B87 : AND3
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N56, A1 => UQVN_N55, A2 => TI4);
UQVB_B88 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N56, A1 => UQVN_N54, A2 => D4);
UQVB_B89 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => TG);
UQVB_B90 : PW
	PORT MAP (PULSE => TG);
UQVB_B91 : SHFE
	PORT MAP (REF => TG, DATA => TI4);
UQVB_B92 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B93 : AND2
	PORT MAP (Z0 => UQVN_N59, A0 => D7, A1 => G);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N63, A0 => G);
UQVB_B95 : PW
	PORT MAP (PULSE => G);
UQVB_B96 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N64);
UQVB_B97 : OR5
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N58, A1 => UQVN_N61, A2 => UQVN_N57, 
	A3 => UQVN_N60, A4 => UQVN_N59);
UQVB_B98 : AND2
	PORT MAP (Z0 => UQVN_N60, A0 => TI7, A1 => TG);
UQVB_B99 : AND3
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N64, A1 => UQVN_N63, A2 => UQVN_N62);
UQVB_B100 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N64, A1 => UQVN_N63, A2 => TI7);
UQVB_B101 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N64, A1 => UQVN_N62, A2 => D7);
UQVB_B102 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => TG);
UQVB_B103 : PW
	PORT MAP (PULSE => TG);
UQVB_B104 : SHFE
	PORT MAP (REF => TG, DATA => TI7);
END lattice_arch;
-- VHDL netlist for LD71
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD71 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        G : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic
    );
END LD71;


ARCHITECTURE lattice_arch OF LD71 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => UQVN_N4, A2 => G);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B4 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B5 : PW
	PORT MAP (PULSE => G);
UQVB_B6 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N9);
UQVB_B9 : OR5
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N7, A4 => UQVN_N3);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N4, A1 => TI0, A2 => TG);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => UQVN_N8);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => TI0);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N8, 
	A3 => D0);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => TG);
UQVB_B15 : PW
	PORT MAP (PULSE => TG);
UQVB_B16 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B17 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD74
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD74 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        G : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD74;


ARCHITECTURE lattice_arch OF LD74 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => UQVN_N4, A2 => G);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B4 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B5 : PW
	PORT MAP (PULSE => G);
UQVB_B6 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N9);
UQVB_B9 : OR5
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N7, A4 => UQVN_N3);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N4, A1 => TI3, A2 => TG);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => UQVN_N8);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => TI3);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N8, 
	A3 => D3);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => TG);
UQVB_B15 : PW
	PORT MAP (PULSE => TG);
UQVB_B16 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B17 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => TG);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => D2, A1 => UQVN_N13, A2 => G);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => CD);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B21 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B22 : PW
	PORT MAP (PULSE => G);
UQVB_B23 : SHFE
	PORT MAP (REF => UQVN_N13, DATA => G);
UQVB_B24 : PW
	PORT MAP (PULSE => UQVN_N13);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N18);
UQVB_B26 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N11, A1 => UQVN_N15, A2 => UQVN_N10, 
	A3 => UQVN_N16, A4 => UQVN_N12);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N13, A1 => TI2, A2 => TG);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N18, A1 => UQVN_N13, A2 => UQVN_N14, 
	A3 => UQVN_N17);
UQVB_B29 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N18, A1 => UQVN_N13, A2 => UQVN_N14, 
	A3 => TI2);
UQVB_B30 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N18, A1 => UQVN_N13, A2 => UQVN_N17, 
	A3 => D2);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TG);
UQVB_B32 : PW
	PORT MAP (PULSE => TG);
UQVB_B33 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B34 : SHFE
	PORT MAP (REF => UQVN_N13, DATA => TG);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D1, A1 => UQVN_N22, A2 => G);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B38 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B39 : PW
	PORT MAP (PULSE => G);
UQVB_B40 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B41 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B42 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N27);
UQVB_B43 : OR5
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N20, A1 => UQVN_N24, A2 => UQVN_N19, 
	A3 => UQVN_N25, A4 => UQVN_N21);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N22, A1 => TI1, A2 => TG);
UQVB_B45 : AND4
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N27, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => UQVN_N26);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N27, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => TI1);
UQVB_B47 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N27, A1 => UQVN_N22, A2 => UQVN_N26, 
	A3 => D1);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => TG);
UQVB_B49 : PW
	PORT MAP (PULSE => TG);
UQVB_B50 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B51 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => TG);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => D0, A1 => UQVN_N31, A2 => G);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => CD);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => G);
UQVB_B55 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B56 : PW
	PORT MAP (PULSE => G);
UQVB_B57 : SHFE
	PORT MAP (REF => UQVN_N31, DATA => G);
UQVB_B58 : PW
	PORT MAP (PULSE => UQVN_N31);
UQVB_B59 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N36);
UQVB_B60 : OR5
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N29, A1 => UQVN_N33, A2 => UQVN_N28, 
	A3 => UQVN_N34, A4 => UQVN_N30);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N31, A1 => TI0, A2 => TG);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N36, A1 => UQVN_N31, A2 => UQVN_N32, 
	A3 => UQVN_N35);
UQVB_B63 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N36, A1 => UQVN_N31, A2 => UQVN_N32, 
	A3 => TI0);
UQVB_B64 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N36, A1 => UQVN_N31, A2 => UQVN_N35, 
	A3 => D0);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => TG);
UQVB_B66 : PW
	PORT MAP (PULSE => TG);
UQVB_B67 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B68 : SHFE
	PORT MAP (REF => UQVN_N31, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD78
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD78 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        G : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD78;


ARCHITECTURE lattice_arch OF LD78 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72 : std_logic;


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => D3, A1 => UQVN_N4, A2 => G);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => CD);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => G);
UQVB_B4 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B5 : PW
	PORT MAP (PULSE => G);
UQVB_B6 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => G);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N4);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N9);
UQVB_B9 : OR5
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N7, A4 => UQVN_N3);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N4, A1 => TI3, A2 => TG);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => UQVN_N8);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => TI3);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N9, A1 => UQVN_N4, A2 => UQVN_N8, 
	A3 => D3);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => TG);
UQVB_B15 : PW
	PORT MAP (PULSE => TG);
UQVB_B16 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B17 : SHFE
	PORT MAP (REF => UQVN_N4, DATA => TG);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => D2, A1 => UQVN_N13, A2 => G);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => CD);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B21 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B22 : PW
	PORT MAP (PULSE => G);
UQVB_B23 : SHFE
	PORT MAP (REF => UQVN_N13, DATA => G);
UQVB_B24 : PW
	PORT MAP (PULSE => UQVN_N13);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N18);
UQVB_B26 : OR5
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N11, A1 => UQVN_N15, A2 => UQVN_N10, 
	A3 => UQVN_N16, A4 => UQVN_N12);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N13, A1 => TI2, A2 => TG);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N18, A1 => UQVN_N13, A2 => UQVN_N14, 
	A3 => UQVN_N17);
UQVB_B29 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N18, A1 => UQVN_N13, A2 => UQVN_N14, 
	A3 => TI2);
UQVB_B30 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N18, A1 => UQVN_N13, A2 => UQVN_N17, 
	A3 => D2);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TG);
UQVB_B32 : PW
	PORT MAP (PULSE => TG);
UQVB_B33 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B34 : SHFE
	PORT MAP (REF => UQVN_N13, DATA => TG);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D1, A1 => UQVN_N22, A2 => G);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => G);
UQVB_B38 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B39 : PW
	PORT MAP (PULSE => G);
UQVB_B40 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B41 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B42 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N27);
UQVB_B43 : OR5
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N20, A1 => UQVN_N24, A2 => UQVN_N19, 
	A3 => UQVN_N25, A4 => UQVN_N21);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N22, A1 => TI1, A2 => TG);
UQVB_B45 : AND4
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N27, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => UQVN_N26);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N27, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => TI1);
UQVB_B47 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N27, A1 => UQVN_N22, A2 => UQVN_N26, 
	A3 => D1);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => TG);
UQVB_B49 : PW
	PORT MAP (PULSE => TG);
UQVB_B50 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B51 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => TG);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => D0, A1 => UQVN_N31, A2 => G);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => CD);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => G);
UQVB_B55 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B56 : PW
	PORT MAP (PULSE => G);
UQVB_B57 : SHFE
	PORT MAP (REF => UQVN_N31, DATA => G);
UQVB_B58 : PW
	PORT MAP (PULSE => UQVN_N31);
UQVB_B59 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N36);
UQVB_B60 : OR5
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N29, A1 => UQVN_N33, A2 => UQVN_N28, 
	A3 => UQVN_N34, A4 => UQVN_N30);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N31, A1 => TI0, A2 => TG);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N36, A1 => UQVN_N31, A2 => UQVN_N32, 
	A3 => UQVN_N35);
UQVB_B63 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N36, A1 => UQVN_N31, A2 => UQVN_N32, 
	A3 => TI0);
UQVB_B64 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N36, A1 => UQVN_N31, A2 => UQVN_N35, 
	A3 => D0);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => TG);
UQVB_B66 : PW
	PORT MAP (PULSE => TG);
UQVB_B67 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B68 : SHFE
	PORT MAP (REF => UQVN_N31, DATA => TG);
UQVB_B69 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => D6, A1 => UQVN_N40, A2 => G);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CD);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => G);
UQVB_B72 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B73 : PW
	PORT MAP (PULSE => G);
UQVB_B74 : SHFE
	PORT MAP (REF => UQVN_N40, DATA => G);
UQVB_B75 : PW
	PORT MAP (PULSE => UQVN_N40);
UQVB_B76 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N45);
UQVB_B77 : OR5
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N38, A1 => UQVN_N42, A2 => UQVN_N37, 
	A3 => UQVN_N43, A4 => UQVN_N39);
UQVB_B78 : AND3
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N40, A1 => TI6, A2 => TG);
UQVB_B79 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N45, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => UQVN_N44);
UQVB_B80 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N45, A1 => UQVN_N40, A2 => UQVN_N41, 
	A3 => TI6);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N45, A1 => UQVN_N40, A2 => UQVN_N44, 
	A3 => D6);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => TG);
UQVB_B83 : PW
	PORT MAP (PULSE => TG);
UQVB_B84 : SHFE
	PORT MAP (REF => TG, DATA => TI6);
UQVB_B85 : SHFE
	PORT MAP (REF => UQVN_N40, DATA => TG);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N48, A0 => D5, A1 => UQVN_N49, A2 => G);
UQVB_B87 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => CD);
UQVB_B88 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => G);
UQVB_B89 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B90 : PW
	PORT MAP (PULSE => G);
UQVB_B91 : SHFE
	PORT MAP (REF => UQVN_N49, DATA => G);
UQVB_B92 : PW
	PORT MAP (PULSE => UQVN_N49);
UQVB_B93 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N54);
UQVB_B94 : OR5
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N47, A1 => UQVN_N51, A2 => UQVN_N46, 
	A3 => UQVN_N52, A4 => UQVN_N48);
UQVB_B95 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N49, A1 => TI5, A2 => TG);
UQVB_B96 : AND4
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N54, A1 => UQVN_N49, A2 => UQVN_N50, 
	A3 => UQVN_N53);
UQVB_B97 : AND4
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N54, A1 => UQVN_N49, A2 => UQVN_N50, 
	A3 => TI5);
UQVB_B98 : AND4
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N54, A1 => UQVN_N49, A2 => UQVN_N53, 
	A3 => D5);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => TG);
UQVB_B100 : PW
	PORT MAP (PULSE => TG);
UQVB_B101 : SHFE
	PORT MAP (REF => TG, DATA => TI5);
UQVB_B102 : SHFE
	PORT MAP (REF => UQVN_N49, DATA => TG);
UQVB_B103 : AND3
	PORT MAP (Z0 => UQVN_N57, A0 => D4, A1 => UQVN_N58, A2 => G);
UQVB_B104 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => CD);
UQVB_B105 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => G);
UQVB_B106 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B107 : PW
	PORT MAP (PULSE => G);
UQVB_B108 : SHFE
	PORT MAP (REF => UQVN_N58, DATA => G);
UQVB_B109 : PW
	PORT MAP (PULSE => UQVN_N58);
UQVB_B110 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N63);
UQVB_B111 : OR5
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N56, A1 => UQVN_N60, A2 => UQVN_N55, 
	A3 => UQVN_N61, A4 => UQVN_N57);
UQVB_B112 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N58, A1 => TI4, A2 => TG);
UQVB_B113 : AND4
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N63, A1 => UQVN_N58, A2 => UQVN_N59, 
	A3 => UQVN_N62);
UQVB_B114 : AND4
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N63, A1 => UQVN_N58, A2 => UQVN_N59, 
	A3 => TI4);
UQVB_B115 : AND4
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N63, A1 => UQVN_N58, A2 => UQVN_N62, 
	A3 => D4);
UQVB_B116 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => TG);
UQVB_B117 : PW
	PORT MAP (PULSE => TG);
UQVB_B118 : SHFE
	PORT MAP (REF => TG, DATA => TI4);
UQVB_B119 : SHFE
	PORT MAP (REF => UQVN_N58, DATA => TG);
UQVB_B120 : AND3
	PORT MAP (Z0 => UQVN_N66, A0 => D7, A1 => UQVN_N67, A2 => G);
UQVB_B121 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => CD);
UQVB_B122 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => G);
UQVB_B123 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B124 : PW
	PORT MAP (PULSE => G);
UQVB_B125 : SHFE
	PORT MAP (REF => UQVN_N67, DATA => G);
UQVB_B126 : PW
	PORT MAP (PULSE => UQVN_N67);
UQVB_B127 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N72);
UQVB_B128 : OR5
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N65, A1 => UQVN_N69, A2 => UQVN_N64, 
	A3 => UQVN_N70, A4 => UQVN_N66);
UQVB_B129 : AND3
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N67, A1 => TI7, A2 => TG);
UQVB_B130 : AND4
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N72, A1 => UQVN_N67, A2 => UQVN_N68, 
	A3 => UQVN_N71);
UQVB_B131 : AND4
	PORT MAP (Z0 => UQVN_N69, A0 => UQVN_N72, A1 => UQVN_N67, A2 => UQVN_N68, 
	A3 => TI7);
UQVB_B132 : AND4
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N72, A1 => UQVN_N67, A2 => UQVN_N71, 
	A3 => D7);
UQVB_B133 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => TG);
UQVB_B134 : PW
	PORT MAP (PULSE => TG);
UQVB_B135 : SHFE
	PORT MAP (REF => TG, DATA => TI7);
UQVB_B136 : SHFE
	PORT MAP (REF => UQVN_N67, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD81
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD81 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic
    );
END LD81;


ARCHITECTURE lattice_arch OF LD81 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D0, A1 => G);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B3 : PW
	PORT MAP (PULSE => G);
UQVB_B4 : PW
	PORT MAP (PULSE => PD);
UQVB_B5 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B6 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N8);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => TI0, A1 => TG);
UQVB_B9 : OR6
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N3, A5 => PD);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N4, A2 => UQVN_N7);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => UQVN_N4, A2 => TI0);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N7, A2 => D0);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => TG);
UQVB_B14 : PW
	PORT MAP (PULSE => TG);
UQVB_B15 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B16 : SHFE
	PORT MAP (REF => PD, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD84
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD84 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD84;


ARCHITECTURE lattice_arch OF LD84 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D2, A1 => G);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B3 : PW
	PORT MAP (PULSE => G);
UQVB_B4 : PW
	PORT MAP (PULSE => PD);
UQVB_B5 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B6 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N8);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => TI2, A1 => TG);
UQVB_B9 : OR6
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N3, A5 => PD);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N4, A2 => UQVN_N7);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => UQVN_N4, A2 => TI2);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N7, A2 => D2);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => TG);
UQVB_B14 : PW
	PORT MAP (PULSE => TG);
UQVB_B15 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B16 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => D3, A1 => G);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => G);
UQVB_B19 : PW
	PORT MAP (PULSE => G);
UQVB_B20 : PW
	PORT MAP (PULSE => PD);
UQVB_B21 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B22 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N16);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => TI3, A1 => TG);
UQVB_B25 : OR6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N10, A1 => UQVN_N9, A2 => UQVN_N14, 
	A3 => UQVN_N13, A4 => UQVN_N11, A5 => PD);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N12, A2 => UQVN_N15);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N16, A1 => UQVN_N12, A2 => TI3);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N16, A1 => UQVN_N15, A2 => D3);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => TG);
UQVB_B30 : PW
	PORT MAP (PULSE => TG);
UQVB_B31 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B32 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D1, A1 => G);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => G);
UQVB_B35 : PW
	PORT MAP (PULSE => G);
UQVB_B36 : PW
	PORT MAP (PULSE => PD);
UQVB_B37 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B38 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B39 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N24);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => TI1, A1 => TG);
UQVB_B41 : OR6
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N22, 
	A3 => UQVN_N21, A4 => UQVN_N19, A5 => PD);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N24, A1 => UQVN_N20, A2 => UQVN_N23);
UQVB_B43 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N24, A1 => UQVN_N20, A2 => TI1);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N24, A1 => UQVN_N23, A2 => D1);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => TG);
UQVB_B46 : PW
	PORT MAP (PULSE => TG);
UQVB_B47 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B48 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B49 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => D0, A1 => G);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => G);
UQVB_B51 : PW
	PORT MAP (PULSE => G);
UQVB_B52 : PW
	PORT MAP (PULSE => PD);
UQVB_B53 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B54 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N32);
UQVB_B56 : AND2
	PORT MAP (Z0 => UQVN_N29, A0 => TI0, A1 => TG);
UQVB_B57 : OR6
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N27, A5 => PD);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N28, A2 => UQVN_N31);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N32, A1 => UQVN_N28, A2 => TI0);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N32, A1 => UQVN_N31, A2 => D0);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => TG);
UQVB_B62 : PW
	PORT MAP (PULSE => TG);
UQVB_B63 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B64 : SHFE
	PORT MAP (REF => PD, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD88
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD88 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD88;


ARCHITECTURE lattice_arch OF LD88 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => D7, A1 => G);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B3 : PW
	PORT MAP (PULSE => G);
UQVB_B4 : PW
	PORT MAP (PULSE => PD);
UQVB_B5 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B6 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N8);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => TI7, A1 => TG);
UQVB_B9 : OR6
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N3, A5 => PD);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => UQVN_N4, A2 => UQVN_N7);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N8, A1 => UQVN_N4, A2 => TI7);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N7, A2 => D7);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => TG);
UQVB_B14 : PW
	PORT MAP (PULSE => TG);
UQVB_B15 : SHFE
	PORT MAP (REF => TG, DATA => TI7);
UQVB_B16 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => D6, A1 => G);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => G);
UQVB_B19 : PW
	PORT MAP (PULSE => G);
UQVB_B20 : PW
	PORT MAP (PULSE => PD);
UQVB_B21 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B22 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B23 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N16);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => TI6, A1 => TG);
UQVB_B25 : OR6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N10, A1 => UQVN_N9, A2 => UQVN_N14, 
	A3 => UQVN_N13, A4 => UQVN_N11, A5 => PD);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N12, A2 => UQVN_N15);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N16, A1 => UQVN_N12, A2 => TI6);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N16, A1 => UQVN_N15, A2 => D6);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => TG);
UQVB_B30 : PW
	PORT MAP (PULSE => TG);
UQVB_B31 : SHFE
	PORT MAP (REF => TG, DATA => TI6);
UQVB_B32 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => D5, A1 => G);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => G);
UQVB_B35 : PW
	PORT MAP (PULSE => G);
UQVB_B36 : PW
	PORT MAP (PULSE => PD);
UQVB_B37 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B38 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B39 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N24);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => TI5, A1 => TG);
UQVB_B41 : OR6
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N22, 
	A3 => UQVN_N21, A4 => UQVN_N19, A5 => PD);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N24, A1 => UQVN_N20, A2 => UQVN_N23);
UQVB_B43 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N24, A1 => UQVN_N20, A2 => TI5);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N24, A1 => UQVN_N23, A2 => D5);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => TG);
UQVB_B46 : PW
	PORT MAP (PULSE => TG);
UQVB_B47 : SHFE
	PORT MAP (REF => TG, DATA => TI5);
UQVB_B48 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B49 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => D4, A1 => G);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => G);
UQVB_B51 : PW
	PORT MAP (PULSE => G);
UQVB_B52 : PW
	PORT MAP (PULSE => PD);
UQVB_B53 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B54 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N32);
UQVB_B56 : AND2
	PORT MAP (Z0 => UQVN_N29, A0 => TI4, A1 => TG);
UQVB_B57 : OR6
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N26, A1 => UQVN_N25, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N27, A5 => PD);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N32, A1 => UQVN_N28, A2 => UQVN_N31);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N32, A1 => UQVN_N28, A2 => TI4);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N32, A1 => UQVN_N31, A2 => D4);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => TG);
UQVB_B62 : PW
	PORT MAP (PULSE => TG);
UQVB_B63 : SHFE
	PORT MAP (REF => TG, DATA => TI4);
UQVB_B64 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B65 : AND2
	PORT MAP (Z0 => UQVN_N35, A0 => D2, A1 => G);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => G);
UQVB_B67 : PW
	PORT MAP (PULSE => G);
UQVB_B68 : PW
	PORT MAP (PULSE => PD);
UQVB_B69 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B70 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B71 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N40);
UQVB_B72 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => TI2, A1 => TG);
UQVB_B73 : OR6
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N34, A1 => UQVN_N33, A2 => UQVN_N38, 
	A3 => UQVN_N37, A4 => UQVN_N35, A5 => PD);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N36, A2 => UQVN_N39);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N36, A2 => TI2);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N40, A1 => UQVN_N39, A2 => D2);
UQVB_B77 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => TG);
UQVB_B78 : PW
	PORT MAP (PULSE => TG);
UQVB_B79 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B80 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B81 : AND2
	PORT MAP (Z0 => UQVN_N43, A0 => D3, A1 => G);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => G);
UQVB_B83 : PW
	PORT MAP (PULSE => G);
UQVB_B84 : PW
	PORT MAP (PULSE => PD);
UQVB_B85 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B86 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B87 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N48);
UQVB_B88 : AND2
	PORT MAP (Z0 => UQVN_N45, A0 => TI3, A1 => TG);
UQVB_B89 : OR6
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N42, A1 => UQVN_N41, A2 => UQVN_N46, 
	A3 => UQVN_N45, A4 => UQVN_N43, A5 => PD);
UQVB_B90 : AND3
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N48, A1 => UQVN_N44, A2 => UQVN_N47);
UQVB_B91 : AND3
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N48, A1 => UQVN_N44, A2 => TI3);
UQVB_B92 : AND3
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N48, A1 => UQVN_N47, A2 => D3);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => TG);
UQVB_B94 : PW
	PORT MAP (PULSE => TG);
UQVB_B95 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B96 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B97 : AND2
	PORT MAP (Z0 => UQVN_N51, A0 => D1, A1 => G);
UQVB_B98 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => G);
UQVB_B99 : PW
	PORT MAP (PULSE => G);
UQVB_B100 : PW
	PORT MAP (PULSE => PD);
UQVB_B101 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B102 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B103 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N56);
UQVB_B104 : AND2
	PORT MAP (Z0 => UQVN_N53, A0 => TI1, A1 => TG);
UQVB_B105 : OR6
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N50, A1 => UQVN_N49, A2 => UQVN_N54, 
	A3 => UQVN_N53, A4 => UQVN_N51, A5 => PD);
UQVB_B106 : AND3
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N56, A1 => UQVN_N52, A2 => UQVN_N55);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N56, A1 => UQVN_N52, A2 => TI1);
UQVB_B108 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N56, A1 => UQVN_N55, A2 => D1);
UQVB_B109 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => TG);
UQVB_B110 : PW
	PORT MAP (PULSE => TG);
UQVB_B111 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B112 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B113 : AND2
	PORT MAP (Z0 => UQVN_N59, A0 => D0, A1 => G);
UQVB_B114 : INV
	PORT MAP (ZN0 => UQVN_N60, A0 => G);
UQVB_B115 : PW
	PORT MAP (PULSE => G);
UQVB_B116 : PW
	PORT MAP (PULSE => PD);
UQVB_B117 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B118 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B119 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N64);
UQVB_B120 : AND2
	PORT MAP (Z0 => UQVN_N61, A0 => TI0, A1 => TG);
UQVB_B121 : OR6
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N58, A1 => UQVN_N57, A2 => UQVN_N62, 
	A3 => UQVN_N61, A4 => UQVN_N59, A5 => PD);
UQVB_B122 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N64, A1 => UQVN_N60, A2 => UQVN_N63);
UQVB_B123 : AND3
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N64, A1 => UQVN_N60, A2 => TI0);
UQVB_B124 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N64, A1 => UQVN_N63, A2 => D0);
UQVB_B125 : INV
	PORT MAP (ZN0 => UQVN_N63, A0 => TG);
UQVB_B126 : PW
	PORT MAP (PULSE => TG);
UQVB_B127 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B128 : SHFE
	PORT MAP (REF => PD, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD91
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD91 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic
    );
END LD91;


ARCHITECTURE lattice_arch OF LD91 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => D0, A1 => UQVN_N2, A2 => G);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N2, A1 => PD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B5 : PW
	PORT MAP (PULSE => G);
UQVB_B6 : PW
	PORT MAP (PULSE => PD);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N2);
UQVB_B8 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => G);
UQVB_B9 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B10 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N10);
UQVB_B12 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => PD);
UQVB_B13 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N1, A5 => UQVN_N3);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => TI0, A1 => UQVN_N2, A2 => TG);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N9);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => TI0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TG);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N9, 
	A3 => D0);
UQVB_B19 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B20 : PW
	PORT MAP (PULSE => TG);
UQVB_B21 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => TG);
UQVB_B22 : SHFE
	PORT MAP (REF => PD, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD94
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD94 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LD94;


ARCHITECTURE lattice_arch OF LD94 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => UQVN_N2, A2 => G);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N2, A1 => PD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B5 : PW
	PORT MAP (PULSE => G);
UQVB_B6 : PW
	PORT MAP (PULSE => PD);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N2);
UQVB_B8 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => G);
UQVB_B9 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B10 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N10);
UQVB_B12 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => PD);
UQVB_B13 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N1, A5 => UQVN_N3);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => TI3, A1 => UQVN_N2, A2 => TG);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N9);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => TI3);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TG);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N9, 
	A3 => D3);
UQVB_B19 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B20 : PW
	PORT MAP (PULSE => TG);
UQVB_B21 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => TG);
UQVB_B22 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CD);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => D2, A1 => UQVN_N12, A2 => G);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N12, A1 => PD);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B27 : PW
	PORT MAP (PULSE => G);
UQVB_B28 : PW
	PORT MAP (PULSE => PD);
UQVB_B29 : PW
	PORT MAP (PULSE => UQVN_N12);
UQVB_B30 : SHFE
	PORT MAP (REF => UQVN_N12, DATA => G);
UQVB_B31 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B32 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N20);
UQVB_B34 : SHFE
	PORT MAP (REF => UQVN_N12, DATA => PD);
UQVB_B35 : OR6
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N16, 
	A3 => UQVN_N15, A4 => UQVN_N11, A5 => UQVN_N13);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => TI2, A1 => UQVN_N12, A2 => TG);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => UQVN_N19);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N20, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => TI2);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => TG);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N12, A2 => UQVN_N19, 
	A3 => D2);
UQVB_B41 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B42 : PW
	PORT MAP (PULSE => TG);
UQVB_B43 : SHFE
	PORT MAP (REF => UQVN_N12, DATA => TG);
UQVB_B44 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D1, A1 => UQVN_N22, A2 => G);
UQVB_B47 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N22, A1 => PD);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => G);
UQVB_B49 : PW
	PORT MAP (PULSE => G);
UQVB_B50 : PW
	PORT MAP (PULSE => PD);
UQVB_B51 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B52 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B53 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B54 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N30);
UQVB_B56 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => PD);
UQVB_B57 : OR6
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N28, A1 => UQVN_N27, A2 => UQVN_N26, 
	A3 => UQVN_N25, A4 => UQVN_N21, A5 => UQVN_N23);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => TI1, A1 => UQVN_N22, A2 => TG);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N30, A1 => UQVN_N22, A2 => UQVN_N24, 
	A3 => UQVN_N29);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N30, A1 => UQVN_N22, A2 => UQVN_N24, 
	A3 => TI1);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => TG);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N30, A1 => UQVN_N22, A2 => UQVN_N29, 
	A3 => D1);
UQVB_B63 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B64 : PW
	PORT MAP (PULSE => TG);
UQVB_B65 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => TG);
UQVB_B66 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => CD);
UQVB_B68 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => D0, A1 => UQVN_N32, A2 => G);
UQVB_B69 : AND2
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N32, A1 => PD);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => G);
UQVB_B71 : PW
	PORT MAP (PULSE => G);
UQVB_B72 : PW
	PORT MAP (PULSE => PD);
UQVB_B73 : PW
	PORT MAP (PULSE => UQVN_N32);
UQVB_B74 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => G);
UQVB_B75 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B76 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B77 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N40);
UQVB_B78 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => PD);
UQVB_B79 : OR6
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35, A4 => UQVN_N31, A5 => UQVN_N33);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => TI0, A1 => UQVN_N32, A2 => TG);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N40, A1 => UQVN_N32, A2 => UQVN_N34, 
	A3 => UQVN_N39);
UQVB_B82 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N40, A1 => UQVN_N32, A2 => UQVN_N34, 
	A3 => TI0);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => TG);
UQVB_B84 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N32, A2 => UQVN_N39, 
	A3 => D0);
UQVB_B85 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B86 : PW
	PORT MAP (PULSE => TG);
UQVB_B87 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => TG);
UQVB_B88 : SHFE
	PORT MAP (REF => PD, DATA => TG);
END lattice_arch;
-- VHDL netlist for LD98
-- Date: 15.5.95 13.46.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LD98 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LD98;


ARCHITECTURE lattice_arch OF LD98 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => UQVN_N2, A2 => G);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N2, A1 => PD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => G);
UQVB_B5 : PW
	PORT MAP (PULSE => G);
UQVB_B6 : PW
	PORT MAP (PULSE => PD);
UQVB_B7 : PW
	PORT MAP (PULSE => UQVN_N2);
UQVB_B8 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => G);
UQVB_B9 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B10 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N10);
UQVB_B12 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => PD);
UQVB_B13 : OR6
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N1, A5 => UQVN_N3);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => TI3, A1 => UQVN_N2, A2 => TG);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N9);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => TI3);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => TG);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N2, A2 => UQVN_N9, 
	A3 => D3);
UQVB_B19 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B20 : PW
	PORT MAP (PULSE => TG);
UQVB_B21 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => TG);
UQVB_B22 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => CD);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => D2, A1 => UQVN_N12, A2 => G);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N12, A1 => PD);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => G);
UQVB_B27 : PW
	PORT MAP (PULSE => G);
UQVB_B28 : PW
	PORT MAP (PULSE => PD);
UQVB_B29 : PW
	PORT MAP (PULSE => UQVN_N12);
UQVB_B30 : SHFE
	PORT MAP (REF => UQVN_N12, DATA => G);
UQVB_B31 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B32 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N20);
UQVB_B34 : SHFE
	PORT MAP (REF => UQVN_N12, DATA => PD);
UQVB_B35 : OR6
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N16, 
	A3 => UQVN_N15, A4 => UQVN_N11, A5 => UQVN_N13);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => TI2, A1 => UQVN_N12, A2 => TG);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => UQVN_N19);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N20, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => TI2);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => TG);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N12, A2 => UQVN_N19, 
	A3 => D2);
UQVB_B41 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B42 : PW
	PORT MAP (PULSE => TG);
UQVB_B43 : SHFE
	PORT MAP (REF => UQVN_N12, DATA => TG);
UQVB_B44 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => CD);
UQVB_B46 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => D1, A1 => UQVN_N22, A2 => G);
UQVB_B47 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N22, A1 => PD);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => G);
UQVB_B49 : PW
	PORT MAP (PULSE => G);
UQVB_B50 : PW
	PORT MAP (PULSE => PD);
UQVB_B51 : PW
	PORT MAP (PULSE => UQVN_N22);
UQVB_B52 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => G);
UQVB_B53 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B54 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B55 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N30);
UQVB_B56 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => PD);
UQVB_B57 : OR6
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N28, A1 => UQVN_N27, A2 => UQVN_N26, 
	A3 => UQVN_N25, A4 => UQVN_N21, A5 => UQVN_N23);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => TI1, A1 => UQVN_N22, A2 => TG);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N30, A1 => UQVN_N22, A2 => UQVN_N24, 
	A3 => UQVN_N29);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N30, A1 => UQVN_N22, A2 => UQVN_N24, 
	A3 => TI1);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => TG);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N30, A1 => UQVN_N22, A2 => UQVN_N29, 
	A3 => D1);
UQVB_B63 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B64 : PW
	PORT MAP (PULSE => TG);
UQVB_B65 : SHFE
	PORT MAP (REF => UQVN_N22, DATA => TG);
UQVB_B66 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => CD);
UQVB_B68 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => D0, A1 => UQVN_N32, A2 => G);
UQVB_B69 : AND2
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N32, A1 => PD);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => G);
UQVB_B71 : PW
	PORT MAP (PULSE => G);
UQVB_B72 : PW
	PORT MAP (PULSE => PD);
UQVB_B73 : PW
	PORT MAP (PULSE => UQVN_N32);
UQVB_B74 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => G);
UQVB_B75 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B76 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B77 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N40);
UQVB_B78 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => PD);
UQVB_B79 : OR6
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35, A4 => UQVN_N31, A5 => UQVN_N33);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => TI0, A1 => UQVN_N32, A2 => TG);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N40, A1 => UQVN_N32, A2 => UQVN_N34, 
	A3 => UQVN_N39);
UQVB_B82 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N40, A1 => UQVN_N32, A2 => UQVN_N34, 
	A3 => TI0);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => TG);
UQVB_B84 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N32, A2 => UQVN_N39, 
	A3 => D0);
UQVB_B85 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B86 : PW
	PORT MAP (PULSE => TG);
UQVB_B87 : SHFE
	PORT MAP (REF => UQVN_N32, DATA => TG);
UQVB_B88 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B89 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => CD);
UQVB_B90 : AND3
	PORT MAP (Z0 => UQVN_N41, A0 => D7, A1 => UQVN_N42, A2 => G);
UQVB_B91 : AND2
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N42, A1 => PD);
UQVB_B92 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => G);
UQVB_B93 : PW
	PORT MAP (PULSE => G);
UQVB_B94 : PW
	PORT MAP (PULSE => PD);
UQVB_B95 : PW
	PORT MAP (PULSE => UQVN_N42);
UQVB_B96 : SHFE
	PORT MAP (REF => UQVN_N42, DATA => G);
UQVB_B97 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B98 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B99 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N50);
UQVB_B100 : SHFE
	PORT MAP (REF => UQVN_N42, DATA => PD);
UQVB_B101 : OR6
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N48, A1 => UQVN_N47, A2 => UQVN_N46, 
	A3 => UQVN_N45, A4 => UQVN_N41, A5 => UQVN_N43);
UQVB_B102 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => TI7, A1 => UQVN_N42, A2 => TG);
UQVB_B103 : AND4
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N50, A1 => UQVN_N42, A2 => UQVN_N44, 
	A3 => UQVN_N49);
UQVB_B104 : AND4
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N50, A1 => UQVN_N42, A2 => UQVN_N44, 
	A3 => TI7);
UQVB_B105 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => TG);
UQVB_B106 : AND4
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N50, A1 => UQVN_N42, A2 => UQVN_N49, 
	A3 => D7);
UQVB_B107 : SHFE
	PORT MAP (REF => TG, DATA => TI7);
UQVB_B108 : PW
	PORT MAP (PULSE => TG);
UQVB_B109 : SHFE
	PORT MAP (REF => UQVN_N42, DATA => TG);
UQVB_B110 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B111 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => CD);
UQVB_B112 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => D6, A1 => UQVN_N52, A2 => G);
UQVB_B113 : AND2
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N52, A1 => PD);
UQVB_B114 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => G);
UQVB_B115 : PW
	PORT MAP (PULSE => G);
UQVB_B116 : PW
	PORT MAP (PULSE => PD);
UQVB_B117 : PW
	PORT MAP (PULSE => UQVN_N52);
UQVB_B118 : SHFE
	PORT MAP (REF => UQVN_N52, DATA => G);
UQVB_B119 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B120 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B121 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N60);
UQVB_B122 : SHFE
	PORT MAP (REF => UQVN_N52, DATA => PD);
UQVB_B123 : OR6
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N58, A1 => UQVN_N57, A2 => UQVN_N56, 
	A3 => UQVN_N55, A4 => UQVN_N51, A5 => UQVN_N53);
UQVB_B124 : AND3
	PORT MAP (Z0 => UQVN_N55, A0 => TI6, A1 => UQVN_N52, A2 => TG);
UQVB_B125 : AND4
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N60, A1 => UQVN_N52, A2 => UQVN_N54, 
	A3 => UQVN_N59);
UQVB_B126 : AND4
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N60, A1 => UQVN_N52, A2 => UQVN_N54, 
	A3 => TI6);
UQVB_B127 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => TG);
UQVB_B128 : AND4
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N60, A1 => UQVN_N52, A2 => UQVN_N59, 
	A3 => D6);
UQVB_B129 : SHFE
	PORT MAP (REF => TG, DATA => TI6);
UQVB_B130 : PW
	PORT MAP (PULSE => TG);
UQVB_B131 : SHFE
	PORT MAP (REF => UQVN_N52, DATA => TG);
UQVB_B132 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B133 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => CD);
UQVB_B134 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => D5, A1 => UQVN_N62, A2 => G);
UQVB_B135 : AND2
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N62, A1 => PD);
UQVB_B136 : INV
	PORT MAP (ZN0 => UQVN_N64, A0 => G);
UQVB_B137 : PW
	PORT MAP (PULSE => G);
UQVB_B138 : PW
	PORT MAP (PULSE => PD);
UQVB_B139 : PW
	PORT MAP (PULSE => UQVN_N62);
UQVB_B140 : SHFE
	PORT MAP (REF => UQVN_N62, DATA => G);
UQVB_B141 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B142 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B143 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N70);
UQVB_B144 : SHFE
	PORT MAP (REF => UQVN_N62, DATA => PD);
UQVB_B145 : OR6
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N68, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => UQVN_N65, A4 => UQVN_N61, A5 => UQVN_N63);
UQVB_B146 : AND3
	PORT MAP (Z0 => UQVN_N65, A0 => TI5, A1 => UQVN_N62, A2 => TG);
UQVB_B147 : AND4
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N70, A1 => UQVN_N62, A2 => UQVN_N64, 
	A3 => UQVN_N69);
UQVB_B148 : AND4
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N70, A1 => UQVN_N62, A2 => UQVN_N64, 
	A3 => TI5);
UQVB_B149 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => TG);
UQVB_B150 : AND4
	PORT MAP (Z0 => UQVN_N68, A0 => UQVN_N70, A1 => UQVN_N62, A2 => UQVN_N69, 
	A3 => D5);
UQVB_B151 : SHFE
	PORT MAP (REF => TG, DATA => TI5);
UQVB_B152 : PW
	PORT MAP (PULSE => TG);
UQVB_B153 : SHFE
	PORT MAP (REF => UQVN_N62, DATA => TG);
UQVB_B154 : SHFE
	PORT MAP (REF => PD, DATA => TG);
UQVB_B155 : INV
	PORT MAP (ZN0 => UQVN_N72, A0 => CD);
UQVB_B156 : AND3
	PORT MAP (Z0 => UQVN_N71, A0 => D4, A1 => UQVN_N72, A2 => G);
UQVB_B157 : AND2
	PORT MAP (Z0 => UQVN_N73, A0 => UQVN_N72, A1 => PD);
UQVB_B158 : INV
	PORT MAP (ZN0 => UQVN_N74, A0 => G);
UQVB_B159 : PW
	PORT MAP (PULSE => G);
UQVB_B160 : PW
	PORT MAP (PULSE => PD);
UQVB_B161 : PW
	PORT MAP (PULSE => UQVN_N72);
UQVB_B162 : SHFE
	PORT MAP (REF => UQVN_N72, DATA => G);
UQVB_B163 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B164 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B165 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N80);
UQVB_B166 : SHFE
	PORT MAP (REF => UQVN_N72, DATA => PD);
UQVB_B167 : OR6
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N78, A1 => UQVN_N77, A2 => UQVN_N76, 
	A3 => UQVN_N75, A4 => UQVN_N71, A5 => UQVN_N73);
UQVB_B168 : AND3
	PORT MAP (Z0 => UQVN_N75, A0 => TI4, A1 => UQVN_N72, A2 => TG);
UQVB_B169 : AND4
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N80, A1 => UQVN_N72, A2 => UQVN_N74, 
	A3 => UQVN_N79);
UQVB_B170 : AND4
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N80, A1 => UQVN_N72, A2 => UQVN_N74, 
	A3 => TI4);
UQVB_B171 : INV
	PORT MAP (ZN0 => UQVN_N79, A0 => TG);
UQVB_B172 : AND4
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N80, A1 => UQVN_N72, A2 => UQVN_N79, 
	A3 => D4);
UQVB_B173 : SHFE
	PORT MAP (REF => TG, DATA => TI4);
UQVB_B174 : PW
	PORT MAP (PULSE => TG);
UQVB_B175 : SHFE
	PORT MAP (REF => UQVN_N72, DATA => TG);
UQVB_B176 : SHFE
	PORT MAP (REF => PD, DATA => TG);
END lattice_arch;
-- VHDL netlist for LDA1
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LDA1 IS 
    PORT (
        D0 : IN std_logic;
        TI0 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic
    );
END LDA1;


ARCHITECTURE lattice_arch OF LDA1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => D0, A1 => UQVN_N2, A2 => G);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => G);
UQVB_B4 : PW
	PORT MAP (PULSE => G);
UQVB_B5 : PW
	PORT MAP (PULSE => PD);
UQVB_B6 : PW
	PORT MAP (PULSE => UQVN_N2);
UQVB_B7 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => G);
UQVB_B8 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B9 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N9);
UQVB_B11 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => PD);
UQVB_B12 : OR6
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N4, A4 => UQVN_N1, A5 => PD);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => TI0, A1 => UQVN_N2, A2 => TG);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N8);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => TI0);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => TG);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N8, 
	A3 => D0);
UQVB_B18 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B19 : PW
	PORT MAP (PULSE => TG);
UQVB_B20 : SHFE
	PORT MAP (REF => PD, DATA => TI0);
UQVB_B21 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => TI0);
END lattice_arch;
-- VHDL netlist for LDA4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LDA4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END LDA4;


ARCHITECTURE lattice_arch OF LDA4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => UQVN_N2, A2 => G);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => G);
UQVB_B4 : PW
	PORT MAP (PULSE => G);
UQVB_B5 : PW
	PORT MAP (PULSE => PD);
UQVB_B6 : PW
	PORT MAP (PULSE => UQVN_N2);
UQVB_B7 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => G);
UQVB_B8 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B9 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N9);
UQVB_B11 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => PD);
UQVB_B12 : OR6
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N4, A4 => UQVN_N1, A5 => PD);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => UQVN_N2, A2 => TG);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N8);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => TI3);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => TG);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N8, 
	A3 => D3);
UQVB_B18 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B19 : PW
	PORT MAP (PULSE => TG);
UQVB_B20 : SHFE
	PORT MAP (REF => PD, DATA => TI3);
UQVB_B21 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => TI3);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => CD);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D2, A1 => UQVN_N11, A2 => G);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => G);
UQVB_B25 : PW
	PORT MAP (PULSE => G);
UQVB_B26 : PW
	PORT MAP (PULSE => PD);
UQVB_B27 : PW
	PORT MAP (PULSE => UQVN_N11);
UQVB_B28 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => G);
UQVB_B29 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B30 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N18);
UQVB_B32 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => PD);
UQVB_B33 : OR6
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N16, A1 => UQVN_N15, A2 => UQVN_N14, 
	A3 => UQVN_N13, A4 => UQVN_N10, A5 => PD);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => TI2, A1 => UQVN_N11, A2 => TG);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N18, A1 => UQVN_N11, A2 => UQVN_N12, 
	A3 => UQVN_N17);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N18, A1 => UQVN_N11, A2 => UQVN_N12, 
	A3 => TI2);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TG);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N18, A1 => UQVN_N11, A2 => UQVN_N17, 
	A3 => D2);
UQVB_B39 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B40 : PW
	PORT MAP (PULSE => TG);
UQVB_B41 : SHFE
	PORT MAP (REF => PD, DATA => TI2);
UQVB_B42 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => TI2);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => CD);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => D1, A1 => UQVN_N20, A2 => G);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => G);
UQVB_B46 : PW
	PORT MAP (PULSE => G);
UQVB_B47 : PW
	PORT MAP (PULSE => PD);
UQVB_B48 : PW
	PORT MAP (PULSE => UQVN_N20);
UQVB_B49 : SHFE
	PORT MAP (REF => UQVN_N20, DATA => G);
UQVB_B50 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B51 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B52 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N27);
UQVB_B53 : SHFE
	PORT MAP (REF => UQVN_N20, DATA => PD);
UQVB_B54 : OR6
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N22, A4 => UQVN_N19, A5 => PD);
UQVB_B55 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => TI1, A1 => UQVN_N20, A2 => TG);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N27, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N26);
UQVB_B57 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N27, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => TI1);
UQVB_B58 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => TG);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N27, A1 => UQVN_N20, A2 => UQVN_N26, 
	A3 => D1);
UQVB_B60 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B61 : PW
	PORT MAP (PULSE => TG);
UQVB_B62 : SHFE
	PORT MAP (REF => PD, DATA => TI1);
UQVB_B63 : SHFE
	PORT MAP (REF => UQVN_N20, DATA => TI1);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => CD);
UQVB_B65 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => D0, A1 => UQVN_N29, A2 => G);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => G);
UQVB_B67 : PW
	PORT MAP (PULSE => G);
UQVB_B68 : PW
	PORT MAP (PULSE => PD);
UQVB_B69 : PW
	PORT MAP (PULSE => UQVN_N29);
UQVB_B70 : SHFE
	PORT MAP (REF => UQVN_N29, DATA => G);
UQVB_B71 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B72 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B73 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N36);
UQVB_B74 : SHFE
	PORT MAP (REF => UQVN_N29, DATA => PD);
UQVB_B75 : OR6
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N34, A1 => UQVN_N33, A2 => UQVN_N32, 
	A3 => UQVN_N31, A4 => UQVN_N28, A5 => PD);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => TI0, A1 => UQVN_N29, A2 => TG);
UQVB_B77 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => UQVN_N29, A2 => UQVN_N30, 
	A3 => UQVN_N35);
UQVB_B78 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N36, A1 => UQVN_N29, A2 => UQVN_N30, 
	A3 => TI0);
UQVB_B79 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => TG);
UQVB_B80 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N36, A1 => UQVN_N29, A2 => UQVN_N35, 
	A3 => D0);
UQVB_B81 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B82 : PW
	PORT MAP (PULSE => TG);
UQVB_B83 : SHFE
	PORT MAP (REF => PD, DATA => TI0);
UQVB_B84 : SHFE
	PORT MAP (REF => UQVN_N29, DATA => TI0);
END lattice_arch;
-- VHDL netlist for LDA8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LDA8 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        TI0 : IN std_logic;
        TI1 : IN std_logic;
        TI2 : IN std_logic;
        TI3 : IN std_logic;
        TI4 : IN std_logic;
        TI5 : IN std_logic;
        TI6 : IN std_logic;
        TI7 : IN std_logic;
        G : IN std_logic;
        PD : IN std_logic;
        CD : IN std_logic;
        TG : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END LDA8;


ARCHITECTURE lattice_arch OF LDA8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT PW
    PORT (
        PULSE : IN std_logic
    );
  END COMPONENT;

for all: PW use  entity  lat_vhd.PW(lattice_arch);


  COMPONENT SHFE
    PORT (
        REF : IN std_logic;
        DATA : IN std_logic
    );
  END COMPONENT;

for all: SHFE use  entity  lat_vhd.SHFE(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => D3, A1 => UQVN_N2, A2 => G);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => G);
UQVB_B4 : PW
	PORT MAP (PULSE => G);
UQVB_B5 : PW
	PORT MAP (PULSE => PD);
UQVB_B6 : PW
	PORT MAP (PULSE => UQVN_N2);
UQVB_B7 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => G);
UQVB_B8 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B9 : SHFE
	PORT MAP (REF => G, DATA => D3);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N9);
UQVB_B11 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => PD);
UQVB_B12 : OR6
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N4, A4 => UQVN_N1, A5 => PD);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => TI3, A1 => UQVN_N2, A2 => TG);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N8);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => TI3);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => TG);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N9, A1 => UQVN_N2, A2 => UQVN_N8, 
	A3 => D3);
UQVB_B18 : SHFE
	PORT MAP (REF => TG, DATA => TI3);
UQVB_B19 : PW
	PORT MAP (PULSE => TG);
UQVB_B20 : SHFE
	PORT MAP (REF => PD, DATA => TI3);
UQVB_B21 : SHFE
	PORT MAP (REF => UQVN_N2, DATA => TI3);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => CD);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D2, A1 => UQVN_N11, A2 => G);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => G);
UQVB_B25 : PW
	PORT MAP (PULSE => G);
UQVB_B26 : PW
	PORT MAP (PULSE => PD);
UQVB_B27 : PW
	PORT MAP (PULSE => UQVN_N11);
UQVB_B28 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => G);
UQVB_B29 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B30 : SHFE
	PORT MAP (REF => G, DATA => D2);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N18);
UQVB_B32 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => PD);
UQVB_B33 : OR6
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N16, A1 => UQVN_N15, A2 => UQVN_N14, 
	A3 => UQVN_N13, A4 => UQVN_N10, A5 => PD);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => TI2, A1 => UQVN_N11, A2 => TG);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N18, A1 => UQVN_N11, A2 => UQVN_N12, 
	A3 => UQVN_N17);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N18, A1 => UQVN_N11, A2 => UQVN_N12, 
	A3 => TI2);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => TG);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N18, A1 => UQVN_N11, A2 => UQVN_N17, 
	A3 => D2);
UQVB_B39 : SHFE
	PORT MAP (REF => TG, DATA => TI2);
UQVB_B40 : PW
	PORT MAP (PULSE => TG);
UQVB_B41 : SHFE
	PORT MAP (REF => PD, DATA => TI2);
UQVB_B42 : SHFE
	PORT MAP (REF => UQVN_N11, DATA => TI2);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => CD);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => D1, A1 => UQVN_N20, A2 => G);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => G);
UQVB_B46 : PW
	PORT MAP (PULSE => G);
UQVB_B47 : PW
	PORT MAP (PULSE => PD);
UQVB_B48 : PW
	PORT MAP (PULSE => UQVN_N20);
UQVB_B49 : SHFE
	PORT MAP (REF => UQVN_N20, DATA => G);
UQVB_B50 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B51 : SHFE
	PORT MAP (REF => G, DATA => D1);
UQVB_B52 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N27);
UQVB_B53 : SHFE
	PORT MAP (REF => UQVN_N20, DATA => PD);
UQVB_B54 : OR6
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N22, A4 => UQVN_N19, A5 => PD);
UQVB_B55 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => TI1, A1 => UQVN_N20, A2 => TG);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N27, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N26);
UQVB_B57 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N27, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => TI1);
UQVB_B58 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => TG);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N27, A1 => UQVN_N20, A2 => UQVN_N26, 
	A3 => D1);
UQVB_B60 : SHFE
	PORT MAP (REF => TG, DATA => TI1);
UQVB_B61 : PW
	PORT MAP (PULSE => TG);
UQVB_B62 : SHFE
	PORT MAP (REF => PD, DATA => TI1);
UQVB_B63 : SHFE
	PORT MAP (REF => UQVN_N20, DATA => TI1);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => CD);
UQVB_B65 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => D0, A1 => UQVN_N29, A2 => G);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => G);
UQVB_B67 : PW
	PORT MAP (PULSE => G);
UQVB_B68 : PW
	PORT MAP (PULSE => PD);
UQVB_B69 : PW
	PORT MAP (PULSE => UQVN_N29);
UQVB_B70 : SHFE
	PORT MAP (REF => UQVN_N29, DATA => G);
UQVB_B71 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B72 : SHFE
	PORT MAP (REF => G, DATA => D0);
UQVB_B73 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N36);
UQVB_B74 : SHFE
	PORT MAP (REF => UQVN_N29, DATA => PD);
UQVB_B75 : OR6
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N34, A1 => UQVN_N33, A2 => UQVN_N32, 
	A3 => UQVN_N31, A4 => UQVN_N28, A5 => PD);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => TI0, A1 => UQVN_N29, A2 => TG);
UQVB_B77 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => UQVN_N29, A2 => UQVN_N30, 
	A3 => UQVN_N35);
UQVB_B78 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N36, A1 => UQVN_N29, A2 => UQVN_N30, 
	A3 => TI0);
UQVB_B79 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => TG);
UQVB_B80 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N36, A1 => UQVN_N29, A2 => UQVN_N35, 
	A3 => D0);
UQVB_B81 : SHFE
	PORT MAP (REF => TG, DATA => TI0);
UQVB_B82 : PW
	PORT MAP (PULSE => TG);
UQVB_B83 : SHFE
	PORT MAP (REF => PD, DATA => TI0);
UQVB_B84 : SHFE
	PORT MAP (REF => UQVN_N29, DATA => TI0);
UQVB_B85 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => CD);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N37, A0 => D7, A1 => UQVN_N38, A2 => G);
UQVB_B87 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => G);
UQVB_B88 : PW
	PORT MAP (PULSE => G);
UQVB_B89 : PW
	PORT MAP (PULSE => PD);
UQVB_B90 : PW
	PORT MAP (PULSE => UQVN_N38);
UQVB_B91 : SHFE
	PORT MAP (REF => UQVN_N38, DATA => G);
UQVB_B92 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B93 : SHFE
	PORT MAP (REF => G, DATA => D7);
UQVB_B94 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N45);
UQVB_B95 : SHFE
	PORT MAP (REF => UQVN_N38, DATA => PD);
UQVB_B96 : OR6
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N43, A1 => UQVN_N42, A2 => UQVN_N41, 
	A3 => UQVN_N40, A4 => UQVN_N37, A5 => PD);
UQVB_B97 : AND3
	PORT MAP (Z0 => UQVN_N40, A0 => TI7, A1 => UQVN_N38, A2 => TG);
UQVB_B98 : AND4
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N45, A1 => UQVN_N38, A2 => UQVN_N39, 
	A3 => UQVN_N44);
UQVB_B99 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N45, A1 => UQVN_N38, A2 => UQVN_N39, 
	A3 => TI7);
UQVB_B100 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => TG);
UQVB_B101 : AND4
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N45, A1 => UQVN_N38, A2 => UQVN_N44, 
	A3 => D7);
UQVB_B102 : SHFE
	PORT MAP (REF => TG, DATA => TI7);
UQVB_B103 : PW
	PORT MAP (PULSE => TG);
UQVB_B104 : SHFE
	PORT MAP (REF => PD, DATA => TI7);
UQVB_B105 : SHFE
	PORT MAP (REF => UQVN_N38, DATA => TI7);
UQVB_B106 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => CD);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N46, A0 => D6, A1 => UQVN_N47, A2 => G);
UQVB_B108 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => G);
UQVB_B109 : PW
	PORT MAP (PULSE => G);
UQVB_B110 : PW
	PORT MAP (PULSE => PD);
UQVB_B111 : PW
	PORT MAP (PULSE => UQVN_N47);
UQVB_B112 : SHFE
	PORT MAP (REF => UQVN_N47, DATA => G);
UQVB_B113 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B114 : SHFE
	PORT MAP (REF => G, DATA => D6);
UQVB_B115 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N54);
UQVB_B116 : SHFE
	PORT MAP (REF => UQVN_N47, DATA => PD);
UQVB_B117 : OR6
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N52, A1 => UQVN_N51, A2 => UQVN_N50, 
	A3 => UQVN_N49, A4 => UQVN_N46, A5 => PD);
UQVB_B118 : AND3
	PORT MAP (Z0 => UQVN_N49, A0 => TI6, A1 => UQVN_N47, A2 => TG);
UQVB_B119 : AND4
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N54, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => UQVN_N53);
UQVB_B120 : AND4
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N54, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => TI6);
UQVB_B121 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => TG);
UQVB_B122 : AND4
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N54, A1 => UQVN_N47, A2 => UQVN_N53, 
	A3 => D6);
UQVB_B123 : SHFE
	PORT MAP (REF => TG, DATA => TI6);
UQVB_B124 : PW
	PORT MAP (PULSE => TG);
UQVB_B125 : SHFE
	PORT MAP (REF => PD, DATA => TI6);
UQVB_B126 : SHFE
	PORT MAP (REF => UQVN_N47, DATA => TI6);
UQVB_B127 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => CD);
UQVB_B128 : AND3
	PORT MAP (Z0 => UQVN_N55, A0 => D5, A1 => UQVN_N56, A2 => G);
UQVB_B129 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => G);
UQVB_B130 : PW
	PORT MAP (PULSE => G);
UQVB_B131 : PW
	PORT MAP (PULSE => PD);
UQVB_B132 : PW
	PORT MAP (PULSE => UQVN_N56);
UQVB_B133 : SHFE
	PORT MAP (REF => UQVN_N56, DATA => G);
UQVB_B134 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B135 : SHFE
	PORT MAP (REF => G, DATA => D5);
UQVB_B136 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N63);
UQVB_B137 : SHFE
	PORT MAP (REF => UQVN_N56, DATA => PD);
UQVB_B138 : OR6
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N61, A1 => UQVN_N60, A2 => UQVN_N59, 
	A3 => UQVN_N58, A4 => UQVN_N55, A5 => PD);
UQVB_B139 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => TI5, A1 => UQVN_N56, A2 => TG);
UQVB_B140 : AND4
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N63, A1 => UQVN_N56, A2 => UQVN_N57, 
	A3 => UQVN_N62);
UQVB_B141 : AND4
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N63, A1 => UQVN_N56, A2 => UQVN_N57, 
	A3 => TI5);
UQVB_B142 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => TG);
UQVB_B143 : AND4
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N63, A1 => UQVN_N56, A2 => UQVN_N62, 
	A3 => D5);
UQVB_B144 : SHFE
	PORT MAP (REF => TG, DATA => TI5);
UQVB_B145 : PW
	PORT MAP (PULSE => TG);
UQVB_B146 : SHFE
	PORT MAP (REF => PD, DATA => TI5);
UQVB_B147 : SHFE
	PORT MAP (REF => UQVN_N56, DATA => TI5);
UQVB_B148 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => CD);
UQVB_B149 : AND3
	PORT MAP (Z0 => UQVN_N64, A0 => D4, A1 => UQVN_N65, A2 => G);
UQVB_B150 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => G);
UQVB_B151 : PW
	PORT MAP (PULSE => G);
UQVB_B152 : PW
	PORT MAP (PULSE => PD);
UQVB_B153 : PW
	PORT MAP (PULSE => UQVN_N65);
UQVB_B154 : SHFE
	PORT MAP (REF => UQVN_N65, DATA => G);
UQVB_B155 : SHFE
	PORT MAP (REF => PD, DATA => G);
UQVB_B156 : SHFE
	PORT MAP (REF => G, DATA => D4);
UQVB_B157 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N72);
UQVB_B158 : SHFE
	PORT MAP (REF => UQVN_N65, DATA => PD);
UQVB_B159 : OR6
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N70, A1 => UQVN_N69, A2 => UQVN_N68, 
	A3 => UQVN_N67, A4 => UQVN_N64, A5 => PD);
UQVB_B160 : AND3
	PORT MAP (Z0 => UQVN_N67, A0 => TI4, A1 => UQVN_N65, A2 => TG);
UQVB_B161 : AND4
	PORT MAP (Z0 => UQVN_N68, A0 => UQVN_N72, A1 => UQVN_N65, A2 => UQVN_N66, 
	A3 => UQVN_N71);
UQVB_B162 : AND4
	PORT MAP (Z0 => UQVN_N69, A0 => UQVN_N72, A1 => UQVN_N65, A2 => UQVN_N66, 
	A3 => TI4);
UQVB_B163 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => TG);
UQVB_B164 : AND4
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N72, A1 => UQVN_N65, A2 => UQVN_N71, 
	A3 => D4);
UQVB_B165 : SHFE
	PORT MAP (REF => TG, DATA => TI4);
UQVB_B166 : PW
	PORT MAP (PULSE => TG);
UQVB_B167 : SHFE
	PORT MAP (REF => PD, DATA => TI4);
UQVB_B168 : SHFE
	PORT MAP (REF => UQVN_N65, DATA => TI4);
END lattice_arch;
-- VHDL netlist for LSR1
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LSR1 IS 
    PORT (
        S0 : IN std_logic;
        R0 : IN std_logic;
        Q0 : OUT std_logic
    );
END LSR1;


ARCHITECTURE lattice_arch OF LSR1 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : NAND2
	PORT MAP (ZN0 => UQVN_N2, A0 => S0, A1 => UQVN_N1);
UQVB_B2 : NAND2
	PORT MAP (ZN0 => UQVN_N1, A0 => R0, A1 => UQVN_N2);
UQVB_B3 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
END lattice_arch;
-- VHDL netlist for LSR2
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY LSR2 IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        R0 : IN std_logic;
        R1 : IN std_logic;
        Q0 : OUT std_logic
    );
END LSR2;


ARCHITECTURE lattice_arch OF LSR2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT NAND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NAND2 use  entity  lat_vhd.NAND2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => S0, A1 => S1);
UQVB_B2 : NAND2
	PORT MAP (ZN0 => UQVN_N2, A0 => UQVN_N4, A1 => UQVN_N1);
UQVB_B3 : NAND2
	PORT MAP (ZN0 => UQVN_N1, A0 => UQVN_N3, A1 => UQVN_N2);
UQVB_B4 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N2);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N3, A0 => R0, A1 => R1);
END lattice_arch;
-- VHDL netlist for MAG2
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MAG2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        GTI : IN std_logic;
        EQI : IN std_logic;
        LTI : IN std_logic;
        GT : OUT std_logic;
        EQ : OUT std_logic;
        LT : OUT std_logic
    );
END MAG2;


ARCHITECTURE lattice_arch OF MAG2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => A0);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => A1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => B0);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => B1);
UQVB_B5 : AND7
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N19, 
	A3 => UQVN_N18, A4 => UQVN_N15, A5 => EQI, A6 => UQVN_N14);
UQVB_B6 : AND7
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N17, A1 => A0, A2 => UQVN_N19, 
	A3 => B0, A4 => UQVN_N15, A5 => EQI, A6 => UQVN_N14);
UQVB_B7 : AND7
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => UQVN_N16, A2 => B1, 
	A3 => UQVN_N18, A4 => UQVN_N15, A5 => EQI, A6 => UQVN_N14);
UQVB_B8 : AND7
	PORT MAP (Z0 => UQVN_N3, A0 => A1, A1 => A0, A2 => B1, 
	A3 => B0, A4 => UQVN_N15, A5 => EQI, A6 => UQVN_N14);
UQVB_B9 : OR4
	PORT MAP (Z0 => EQ, A0 => UQVN_N4, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N15, A1 => UQVN_N13, A2 => GTI);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => LTI, A1 => UQVN_N13, A2 => UQVN_N14);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N17, A1 => UQVN_N16, A2 => B0, 
	A3 => UQVN_N15, A4 => EQI, A5 => UQVN_N14);
UQVB_B13 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N16, A1 => B1, A2 => B0, 
	A3 => UQVN_N15, A4 => EQI, A5 => UQVN_N14);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => GTI);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => EQI);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => LTI);
UQVB_B17 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => A1, A1 => UQVN_N19, A2 => UQVN_N15, 
	A3 => EQI, A4 => UQVN_N14);
UQVB_B18 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => UQVN_N19, A2 => UQVN_N18, 
	A3 => UQVN_N15, A4 => EQI, A5 => UQVN_N14);
UQVB_B19 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => A1, A1 => A0, A2 => UQVN_N18, 
	A3 => UQVN_N15, A4 => EQI, A5 => UQVN_N14);
UQVB_B20 : OR4
	PORT MAP (Z0 => GT, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N8);
UQVB_B21 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N17, A1 => B1, A2 => UQVN_N15, 
	A3 => EQI, A4 => UQVN_N14);
UQVB_B22 : OR4
	PORT MAP (Z0 => LT, A0 => UQVN_N9, A1 => UQVN_N10, A2 => UQVN_N12, 
	A3 => UQVN_N11);
END lattice_arch;
-- VHDL netlist for MAG4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MAG4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        GTI : IN std_logic;
        EQI : IN std_logic;
        LTI : IN std_logic;
        GT : OUT std_logic;
        EQ : OUT std_logic;
        LT : OUT std_logic
    );
END MAG4;


ARCHITECTURE lattice_arch OF MAG4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LTI);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => GTI);
UQVB_B3 : AND11
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B4 : AND11
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => A0, A4 => UQVN_N73, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B5 : AND11
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N69, A1 => UQVN_N68, A2 => A1, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => UQVN_N72, A6 => B1, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B6 : AND11
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N69, A1 => UQVN_N68, A2 => A1, 
	A3 => A0, A4 => UQVN_N73, A5 => UQVN_N72, A6 => B1, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B7 : AND11
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N69, A1 => A2, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => B2, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B8 : AND11
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N69, A1 => A2, A2 => UQVN_N67, 
	A3 => A0, A4 => UQVN_N73, A5 => B2, A6 => UQVN_N71, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B9 : AND11
	PORT MAP (Z0 => UQVN_N9, A0 => A3, A1 => UQVN_N68, A2 => A1, 
	A3 => A0, A4 => B3, A5 => UQVN_N72, A6 => B1, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B10 : AND11
	PORT MAP (Z0 => UQVN_N10, A0 => A3, A1 => UQVN_N68, A2 => A1, 
	A3 => UQVN_N66, A4 => B3, A5 => UQVN_N72, A6 => B1, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B11 : AND11
	PORT MAP (Z0 => UQVN_N11, A0 => A3, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => A0, A4 => B3, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B12 : AND11
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N69, A1 => A2, A2 => A1, 
	A3 => A0, A4 => UQVN_N73, A5 => B2, A6 => B1, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B13 : AND11
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N69, A1 => A2, A2 => A1, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => B2, A6 => B1, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B14 : AND11
	PORT MAP (Z0 => UQVN_N12, A0 => A3, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => B3, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B15 : AND11
	PORT MAP (Z0 => UQVN_N21, A0 => A3, A1 => A2, A2 => A1, 
	A3 => A0, A4 => B3, A5 => B2, A6 => B1, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B16 : AND11
	PORT MAP (Z0 => UQVN_N17, A0 => A3, A1 => A2, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => B3, A5 => B2, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B17 : AND11
	PORT MAP (Z0 => UQVN_N16, A0 => A3, A1 => A2, A2 => UQVN_N67, 
	A3 => A0, A4 => B3, A5 => B2, A6 => UQVN_N71, 
	A7 => B0, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B18 : AND11
	PORT MAP (Z0 => UQVN_N15, A0 => A3, A1 => A2, A2 => A1, 
	A3 => UQVN_N66, A4 => B3, A5 => B2, A6 => B1, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B19 : OR7
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N9, A1 => UQVN_N5, A2 => UQVN_N4, 
	A3 => UQVN_N3, A4 => UQVN_N6, A5 => UQVN_N7, A6 => UQVN_N8);
UQVB_B20 : OR5
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N10);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N15, 
	A3 => UQVN_N21);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N73, A0 => B3);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N72, A0 => B2);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => B1);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => B0);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => A1);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => A0);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => A2);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => A3);
UQVB_B30 : OR3
	PORT MAP (Z0 => EQ, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B31 : AND7
	PORT MAP (Z0 => UQVN_N32, A0 => A2, A1 => A1, A2 => UQVN_N73, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B32 : AND7
	PORT MAP (Z0 => UQVN_N30, A0 => A3, A1 => A1, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B33 : AND7
	PORT MAP (Z0 => UQVN_N31, A0 => A3, A1 => A2, A2 => A1, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B34 : AND6
	PORT MAP (Z0 => UQVN_N37, A0 => A2, A1 => UQVN_N73, A2 => UQVN_N72, 
	A3 => UQVN_N43, A4 => EQI, A5 => UQVN_N42);
UQVB_B35 : AND6
	PORT MAP (Z0 => UQVN_N36, A0 => A3, A1 => A2, A2 => UQVN_N72, 
	A3 => UQVN_N43, A4 => EQI, A5 => UQVN_N42);
UQVB_B36 : AND5
	PORT MAP (Z0 => UQVN_N35, A0 => A3, A1 => UQVN_N73, A2 => UQVN_N43, 
	A3 => EQI, A4 => UQVN_N42);
UQVB_B37 : OR7
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N29, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => UQVN_N24, A5 => UQVN_N22, A6 => UQVN_N23);
UQVB_B38 : OR5
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N34, A1 => UQVN_N33, A2 => UQVN_N32, 
	A3 => UQVN_N30, A4 => UQVN_N31);
UQVB_B39 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => GTI, A1 => UQVN_N25, A2 => UQVN_N43);
UQVB_B40 : OR4
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => LTI);
UQVB_B42 : OR3
	PORT MAP (Z0 => GT, A0 => UQVN_N41, A1 => UQVN_N39, A2 => UQVN_N40);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => EQI);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => GTI);
UQVB_B45 : AND8
	PORT MAP (Z0 => UQVN_N29, A0 => A0, A1 => UQVN_N73, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B46 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => A1, A1 => A0, A2 => UQVN_N73, 
	A3 => UQVN_N72, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B47 : AND8
	PORT MAP (Z0 => UQVN_N27, A0 => A2, A1 => A0, A2 => UQVN_N73, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B48 : AND8
	PORT MAP (Z0 => UQVN_N26, A0 => A3, A1 => A0, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B49 : AND8
	PORT MAP (Z0 => UQVN_N24, A0 => A2, A1 => A1, A2 => A0, 
	A3 => UQVN_N73, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B50 : AND8
	PORT MAP (Z0 => UQVN_N22, A0 => A3, A1 => A1, A2 => A0, 
	A3 => UQVN_N72, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B51 : AND8
	PORT MAP (Z0 => UQVN_N23, A0 => A3, A1 => A2, A2 => A0, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B52 : AND7
	PORT MAP (Z0 => UQVN_N33, A0 => A1, A1 => UQVN_N73, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B53 : AND8
	PORT MAP (Z0 => UQVN_N34, A0 => A3, A1 => A2, A2 => A1, 
	A3 => A0, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B54 : AND8
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N69, A1 => UQVN_N66, A2 => B2, 
	A3 => B1, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B55 : AND8
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N68, A1 => UQVN_N66, A2 => B3, 
	A3 => B1, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B56 : AND8
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N67, A1 => UQVN_N66, A2 => B3, 
	A3 => B2, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B57 : AND8
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N66, A1 => B3, A2 => B2, 
	A3 => B1, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B58 : AND7
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => B1, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B59 : AND7
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N69, A1 => UQVN_N67, A2 => B2, 
	A3 => B1, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B60 : AND7
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N68, A1 => UQVN_N67, A2 => B3, 
	A3 => B1, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B61 : AND7
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N67, A1 => B3, A2 => B2, 
	A3 => B1, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B62 : OR7
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N46, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => UQVN_N49, A4 => UQVN_N50, A5 => UQVN_N51, A6 => UQVN_N52);
UQVB_B63 : OR5
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N53, A1 => UQVN_N54, A2 => UQVN_N55, 
	A3 => UQVN_N56, A4 => UQVN_N57);
UQVB_B64 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N44, A1 => UQVN_N65, A2 => LTI);
UQVB_B65 : AND6
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N69, A1 => UQVN_N68, A2 => B2, 
	A3 => UQVN_N45, A4 => EQI, A5 => UQVN_N44);
UQVB_B66 : AND6
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N68, A1 => B3, A2 => B2, 
	A3 => UQVN_N45, A4 => EQI, A5 => UQVN_N44);
UQVB_B67 : AND5
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N69, A1 => B3, A2 => UQVN_N45, 
	A3 => EQI, A4 => UQVN_N44);
UQVB_B68 : OR4
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N61, A1 => UQVN_N60, A2 => UQVN_N59, 
	A3 => UQVN_N58);
UQVB_B69 : OR3
	PORT MAP (Z0 => LT, A0 => UQVN_N63, A1 => UQVN_N62, A2 => UQVN_N64);
UQVB_B70 : AND8
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => LTI);
UQVB_B72 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => EQI);
UQVB_B73 : AND8
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N66, 
	A3 => B1, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B74 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => GTI);
UQVB_B75 : AND8
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N69, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => B2, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B76 : AND8
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N68, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => B3, A4 => B0, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
END lattice_arch;
-- VHDL netlist for MAG8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MAG8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        GTI : IN std_logic;
        EQI : IN std_logic;
        LTI : IN std_logic;
        GT : OUT std_logic;
        EQ : OUT std_logic;
        LT : OUT std_logic
    );
END MAG8;


ARCHITECTURE lattice_arch OF MAG8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 UQVN_N113, UQVN_N114, UQVN_N115, UQVN_N116,
	 UQVN_N117, UQVN_N118, UQVN_N119, UQVN_N120,
	 UQVN_N121, UQVN_N122, UQVN_N123, UQVN_N124,
	 UQVN_N125, UQVN_N126, UQVN_N127, UQVN_N128,
	 UQVN_N129, UQVN_N130, UQVN_N131, UQVN_N132,
	 UQVN_N133, UQVN_N134, UQVN_N135, UQVN_N136,
	 UQVN_N137, UQVN_N138, UQVN_N139, UQVN_N140,
	 UQVN_N141, UQVN_N142, UQVN_N143, UQVN_N144,
	 UQVN_N145, UQVN_N146, UQVN_N147, UQVN_N148,
	 UQVN_N149 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND11
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND11 use  entity  lat_vhd.AND11(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LTI);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => GTI);
UQVB_B3 : AND11
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B4 : AND11
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => A4, A4 => UQVN_N73, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B5 : AND11
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N69, A1 => UQVN_N68, A2 => A5, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => UQVN_N72, A6 => B5, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B6 : AND11
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N69, A1 => UQVN_N68, A2 => A5, 
	A3 => A4, A4 => UQVN_N73, A5 => UQVN_N72, A6 => B5, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B7 : AND11
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N69, A1 => A6, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => B6, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B8 : AND11
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N69, A1 => A6, A2 => UQVN_N67, 
	A3 => A4, A4 => UQVN_N73, A5 => B6, A6 => UQVN_N71, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B9 : AND11
	PORT MAP (Z0 => UQVN_N9, A0 => A7, A1 => UQVN_N68, A2 => A5, 
	A3 => A4, A4 => B7, A5 => UQVN_N72, A6 => B5, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B10 : AND11
	PORT MAP (Z0 => UQVN_N10, A0 => A7, A1 => UQVN_N68, A2 => A5, 
	A3 => UQVN_N66, A4 => B7, A5 => UQVN_N72, A6 => B5, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B11 : AND11
	PORT MAP (Z0 => UQVN_N11, A0 => A7, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => A4, A4 => B7, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B12 : AND11
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N69, A1 => A6, A2 => A5, 
	A3 => A4, A4 => UQVN_N73, A5 => B6, A6 => B5, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B13 : AND11
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N69, A1 => A6, A2 => A5, 
	A3 => UQVN_N66, A4 => UQVN_N73, A5 => B6, A6 => B5, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B14 : AND11
	PORT MAP (Z0 => UQVN_N12, A0 => A7, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => B7, A5 => UQVN_N72, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B15 : AND11
	PORT MAP (Z0 => UQVN_N21, A0 => A7, A1 => A6, A2 => A5, 
	A3 => A4, A4 => B7, A5 => B6, A6 => B5, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B16 : AND11
	PORT MAP (Z0 => UQVN_N17, A0 => A7, A1 => A6, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => B7, A5 => B6, A6 => UQVN_N71, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B17 : AND11
	PORT MAP (Z0 => UQVN_N16, A0 => A7, A1 => A6, A2 => UQVN_N67, 
	A3 => A4, A4 => B7, A5 => B6, A6 => UQVN_N71, 
	A7 => B4, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B18 : AND11
	PORT MAP (Z0 => UQVN_N15, A0 => A7, A1 => A6, A2 => A5, 
	A3 => UQVN_N66, A4 => B7, A5 => B6, A6 => B5, 
	A7 => UQVN_N70, A8 => UQVN_N2, A9 => EQI, A10 => UQVN_N1);
UQVB_B19 : OR7
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N9, A1 => UQVN_N5, A2 => UQVN_N4, 
	A3 => UQVN_N3, A4 => UQVN_N6, A5 => UQVN_N7, A6 => UQVN_N8);
UQVB_B20 : OR5
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N12, 
	A3 => UQVN_N11, A4 => UQVN_N10);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N15, 
	A3 => UQVN_N21);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N73, A0 => B7);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N72, A0 => B6);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => B5);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => B4);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => A5);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => A4);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => A6);
UQVB_B29 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => A7);
UQVB_B30 : OR3
	PORT MAP (Z0 => UQVN_N148, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B31 : AND7
	PORT MAP (Z0 => UQVN_N32, A0 => A6, A1 => A5, A2 => UQVN_N73, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B32 : AND7
	PORT MAP (Z0 => UQVN_N30, A0 => A7, A1 => A5, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B33 : AND7
	PORT MAP (Z0 => UQVN_N31, A0 => A7, A1 => A6, A2 => A5, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B34 : AND6
	PORT MAP (Z0 => UQVN_N37, A0 => A6, A1 => UQVN_N73, A2 => UQVN_N72, 
	A3 => UQVN_N43, A4 => EQI, A5 => UQVN_N42);
UQVB_B35 : AND6
	PORT MAP (Z0 => UQVN_N36, A0 => A7, A1 => A6, A2 => UQVN_N72, 
	A3 => UQVN_N43, A4 => EQI, A5 => UQVN_N42);
UQVB_B36 : AND5
	PORT MAP (Z0 => UQVN_N35, A0 => A7, A1 => UQVN_N73, A2 => UQVN_N43, 
	A3 => EQI, A4 => UQVN_N42);
UQVB_B37 : OR7
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N29, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => UQVN_N24, A5 => UQVN_N22, A6 => UQVN_N23);
UQVB_B38 : OR5
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N34, A1 => UQVN_N33, A2 => UQVN_N32, 
	A3 => UQVN_N30, A4 => UQVN_N31);
UQVB_B39 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => GTI, A1 => UQVN_N25, A2 => UQVN_N43);
UQVB_B40 : OR4
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N36, 
	A3 => UQVN_N35);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => LTI);
UQVB_B42 : OR3
	PORT MAP (Z0 => UQVN_N147, A0 => UQVN_N41, A1 => UQVN_N39, A2 => UQVN_N40);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => EQI);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => GTI);
UQVB_B45 : AND8
	PORT MAP (Z0 => UQVN_N29, A0 => A4, A1 => UQVN_N73, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B46 : AND8
	PORT MAP (Z0 => UQVN_N28, A0 => A5, A1 => A4, A2 => UQVN_N73, 
	A3 => UQVN_N72, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B47 : AND8
	PORT MAP (Z0 => UQVN_N27, A0 => A6, A1 => A4, A2 => UQVN_N73, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B48 : AND8
	PORT MAP (Z0 => UQVN_N26, A0 => A7, A1 => A4, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B49 : AND8
	PORT MAP (Z0 => UQVN_N24, A0 => A6, A1 => A5, A2 => A4, 
	A3 => UQVN_N73, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B50 : AND8
	PORT MAP (Z0 => UQVN_N22, A0 => A7, A1 => A5, A2 => A4, 
	A3 => UQVN_N72, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B51 : AND8
	PORT MAP (Z0 => UQVN_N23, A0 => A7, A1 => A6, A2 => A4, 
	A3 => UQVN_N71, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B52 : AND7
	PORT MAP (Z0 => UQVN_N33, A0 => A5, A1 => UQVN_N73, A2 => UQVN_N72, 
	A3 => UQVN_N71, A4 => UQVN_N43, A5 => EQI, A6 => UQVN_N42);
UQVB_B53 : AND8
	PORT MAP (Z0 => UQVN_N34, A0 => A7, A1 => A6, A2 => A5, 
	A3 => A4, A4 => UQVN_N70, A5 => UQVN_N43, A6 => EQI, 
	A7 => UQVN_N42);
UQVB_B54 : AND8
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N69, A1 => UQVN_N66, A2 => B6, 
	A3 => B5, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B55 : AND8
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N68, A1 => UQVN_N66, A2 => B7, 
	A3 => B5, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B56 : AND8
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N67, A1 => UQVN_N66, A2 => B7, 
	A3 => B6, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B57 : AND8
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N66, A1 => B7, A2 => B6, 
	A3 => B5, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B58 : AND7
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => B5, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B59 : AND7
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N69, A1 => UQVN_N67, A2 => B6, 
	A3 => B5, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B60 : AND7
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N68, A1 => UQVN_N67, A2 => B7, 
	A3 => B5, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B61 : AND7
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N67, A1 => B7, A2 => B6, 
	A3 => B5, A4 => UQVN_N45, A5 => EQI, A6 => UQVN_N44);
UQVB_B62 : OR7
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N46, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => UQVN_N49, A4 => UQVN_N50, A5 => UQVN_N51, A6 => UQVN_N52);
UQVB_B63 : OR5
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N53, A1 => UQVN_N54, A2 => UQVN_N55, 
	A3 => UQVN_N56, A4 => UQVN_N57);
UQVB_B64 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N44, A1 => UQVN_N65, A2 => LTI);
UQVB_B65 : AND6
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N69, A1 => UQVN_N68, A2 => B6, 
	A3 => UQVN_N45, A4 => EQI, A5 => UQVN_N44);
UQVB_B66 : AND6
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N68, A1 => B7, A2 => B6, 
	A3 => UQVN_N45, A4 => EQI, A5 => UQVN_N44);
UQVB_B67 : AND5
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N69, A1 => B7, A2 => UQVN_N45, 
	A3 => EQI, A4 => UQVN_N44);
UQVB_B68 : OR4
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N61, A1 => UQVN_N60, A2 => UQVN_N59, 
	A3 => UQVN_N58);
UQVB_B69 : OR3
	PORT MAP (Z0 => UQVN_N149, A0 => UQVN_N63, A1 => UQVN_N62, A2 => UQVN_N64);
UQVB_B70 : AND8
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N67, 
	A3 => UQVN_N66, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => LTI);
UQVB_B72 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => EQI);
UQVB_B73 : AND8
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N69, A1 => UQVN_N68, A2 => UQVN_N66, 
	A3 => B5, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B74 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => GTI);
UQVB_B75 : AND8
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N69, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => B6, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B76 : AND8
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N68, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => B7, A4 => B4, A5 => UQVN_N45, A6 => EQI, 
	A7 => UQVN_N44);
UQVB_B77 : INV
	PORT MAP (ZN0 => UQVN_N75, A0 => UQVN_N149);
UQVB_B78 : INV
	PORT MAP (ZN0 => UQVN_N74, A0 => UQVN_N147);
UQVB_B79 : AND11
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N142, A1 => UQVN_N141, A2 => UQVN_N140, 
	A3 => UQVN_N139, A4 => UQVN_N146, A5 => UQVN_N145, A6 => UQVN_N144, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B80 : AND11
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N142, A1 => UQVN_N141, A2 => UQVN_N140, 
	A3 => A0, A4 => UQVN_N146, A5 => UQVN_N145, A6 => UQVN_N144, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B81 : AND11
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N142, A1 => UQVN_N141, A2 => A1, 
	A3 => UQVN_N139, A4 => UQVN_N146, A5 => UQVN_N145, A6 => B1, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B82 : AND11
	PORT MAP (Z0 => UQVN_N79, A0 => UQVN_N142, A1 => UQVN_N141, A2 => A1, 
	A3 => A0, A4 => UQVN_N146, A5 => UQVN_N145, A6 => B1, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B83 : AND11
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N142, A1 => A2, A2 => UQVN_N140, 
	A3 => UQVN_N139, A4 => UQVN_N146, A5 => B2, A6 => UQVN_N144, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B84 : AND11
	PORT MAP (Z0 => UQVN_N81, A0 => UQVN_N142, A1 => A2, A2 => UQVN_N140, 
	A3 => A0, A4 => UQVN_N146, A5 => B2, A6 => UQVN_N144, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B85 : AND11
	PORT MAP (Z0 => UQVN_N82, A0 => A3, A1 => UQVN_N141, A2 => A1, 
	A3 => A0, A4 => B3, A5 => UQVN_N145, A6 => B1, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B86 : AND11
	PORT MAP (Z0 => UQVN_N83, A0 => A3, A1 => UQVN_N141, A2 => A1, 
	A3 => UQVN_N139, A4 => B3, A5 => UQVN_N145, A6 => B1, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B87 : AND11
	PORT MAP (Z0 => UQVN_N84, A0 => A3, A1 => UQVN_N141, A2 => UQVN_N140, 
	A3 => A0, A4 => B3, A5 => UQVN_N145, A6 => UQVN_N144, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B88 : AND11
	PORT MAP (Z0 => UQVN_N86, A0 => UQVN_N142, A1 => A2, A2 => A1, 
	A3 => A0, A4 => UQVN_N146, A5 => B2, A6 => B1, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B89 : AND11
	PORT MAP (Z0 => UQVN_N87, A0 => UQVN_N142, A1 => A2, A2 => A1, 
	A3 => UQVN_N139, A4 => UQVN_N146, A5 => B2, A6 => B1, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B90 : AND11
	PORT MAP (Z0 => UQVN_N85, A0 => A3, A1 => UQVN_N141, A2 => UQVN_N140, 
	A3 => UQVN_N139, A4 => B3, A5 => UQVN_N145, A6 => UQVN_N144, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B91 : AND11
	PORT MAP (Z0 => UQVN_N94, A0 => A3, A1 => A2, A2 => A1, 
	A3 => A0, A4 => B3, A5 => B2, A6 => B1, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B92 : AND11
	PORT MAP (Z0 => UQVN_N90, A0 => A3, A1 => A2, A2 => UQVN_N140, 
	A3 => UQVN_N139, A4 => B3, A5 => B2, A6 => UQVN_N144, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B93 : AND11
	PORT MAP (Z0 => UQVN_N89, A0 => A3, A1 => A2, A2 => UQVN_N140, 
	A3 => A0, A4 => B3, A5 => B2, A6 => UQVN_N144, 
	A7 => B0, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B94 : AND11
	PORT MAP (Z0 => UQVN_N88, A0 => A3, A1 => A2, A2 => A1, 
	A3 => UQVN_N139, A4 => B3, A5 => B2, A6 => B1, 
	A7 => UQVN_N143, A8 => UQVN_N75, A9 => UQVN_N148, A10 => UQVN_N74);
UQVB_B95 : OR7
	PORT MAP (Z0 => UQVN_N91, A0 => UQVN_N82, A1 => UQVN_N78, A2 => UQVN_N77, 
	A3 => UQVN_N76, A4 => UQVN_N79, A5 => UQVN_N80, A6 => UQVN_N81);
UQVB_B96 : OR5
	PORT MAP (Z0 => UQVN_N92, A0 => UQVN_N87, A1 => UQVN_N86, A2 => UQVN_N85, 
	A3 => UQVN_N84, A4 => UQVN_N83);
UQVB_B97 : OR4
	PORT MAP (Z0 => UQVN_N93, A0 => UQVN_N90, A1 => UQVN_N89, A2 => UQVN_N88, 
	A3 => UQVN_N94);
UQVB_B98 : INV
	PORT MAP (ZN0 => UQVN_N146, A0 => B3);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N145, A0 => B2);
UQVB_B100 : INV
	PORT MAP (ZN0 => UQVN_N144, A0 => B1);
UQVB_B101 : INV
	PORT MAP (ZN0 => UQVN_N143, A0 => B0);
UQVB_B102 : INV
	PORT MAP (ZN0 => UQVN_N140, A0 => A1);
UQVB_B103 : INV
	PORT MAP (ZN0 => UQVN_N139, A0 => A0);
UQVB_B104 : INV
	PORT MAP (ZN0 => UQVN_N141, A0 => A2);
UQVB_B105 : INV
	PORT MAP (ZN0 => UQVN_N142, A0 => A3);
UQVB_B106 : OR3
	PORT MAP (Z0 => EQ, A0 => UQVN_N93, A1 => UQVN_N92, A2 => UQVN_N91);
UQVB_B107 : AND7
	PORT MAP (Z0 => UQVN_N105, A0 => A2, A1 => A1, A2 => UQVN_N146, 
	A3 => UQVN_N144, A4 => UQVN_N116, A5 => UQVN_N148, A6 => UQVN_N115);
UQVB_B108 : AND7
	PORT MAP (Z0 => UQVN_N103, A0 => A3, A1 => A1, A2 => UQVN_N145, 
	A3 => UQVN_N144, A4 => UQVN_N116, A5 => UQVN_N148, A6 => UQVN_N115);
UQVB_B109 : AND7
	PORT MAP (Z0 => UQVN_N104, A0 => A3, A1 => A2, A2 => A1, 
	A3 => UQVN_N144, A4 => UQVN_N116, A5 => UQVN_N148, A6 => UQVN_N115);
UQVB_B110 : AND6
	PORT MAP (Z0 => UQVN_N110, A0 => A2, A1 => UQVN_N146, A2 => UQVN_N145, 
	A3 => UQVN_N116, A4 => UQVN_N148, A5 => UQVN_N115);
UQVB_B111 : AND6
	PORT MAP (Z0 => UQVN_N109, A0 => A3, A1 => A2, A2 => UQVN_N145, 
	A3 => UQVN_N116, A4 => UQVN_N148, A5 => UQVN_N115);
UQVB_B112 : AND5
	PORT MAP (Z0 => UQVN_N108, A0 => A3, A1 => UQVN_N146, A2 => UQVN_N116, 
	A3 => UQVN_N148, A4 => UQVN_N115);
UQVB_B113 : OR7
	PORT MAP (Z0 => UQVN_N113, A0 => UQVN_N102, A1 => UQVN_N101, A2 => UQVN_N100, 
	A3 => UQVN_N99, A4 => UQVN_N97, A5 => UQVN_N95, A6 => UQVN_N96);
UQVB_B114 : OR5
	PORT MAP (Z0 => UQVN_N112, A0 => UQVN_N107, A1 => UQVN_N106, A2 => UQVN_N105, 
	A3 => UQVN_N103, A4 => UQVN_N104);
UQVB_B115 : AND3
	PORT MAP (Z0 => UQVN_N111, A0 => UQVN_N147, A1 => UQVN_N98, A2 => UQVN_N116);
UQVB_B116 : OR4
	PORT MAP (Z0 => UQVN_N114, A0 => UQVN_N111, A1 => UQVN_N110, A2 => UQVN_N109, 
	A3 => UQVN_N108);
UQVB_B117 : INV
	PORT MAP (ZN0 => UQVN_N116, A0 => UQVN_N149);
UQVB_B118 : OR3
	PORT MAP (Z0 => GT, A0 => UQVN_N114, A1 => UQVN_N112, A2 => UQVN_N113);
UQVB_B119 : INV
	PORT MAP (ZN0 => UQVN_N98, A0 => UQVN_N148);
UQVB_B120 : INV
	PORT MAP (ZN0 => UQVN_N115, A0 => UQVN_N147);
UQVB_B121 : AND8
	PORT MAP (Z0 => UQVN_N102, A0 => A0, A1 => UQVN_N146, A2 => UQVN_N145, 
	A3 => UQVN_N144, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B122 : AND8
	PORT MAP (Z0 => UQVN_N101, A0 => A1, A1 => A0, A2 => UQVN_N146, 
	A3 => UQVN_N145, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B123 : AND8
	PORT MAP (Z0 => UQVN_N100, A0 => A2, A1 => A0, A2 => UQVN_N146, 
	A3 => UQVN_N144, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B124 : AND8
	PORT MAP (Z0 => UQVN_N99, A0 => A3, A1 => A0, A2 => UQVN_N145, 
	A3 => UQVN_N144, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B125 : AND8
	PORT MAP (Z0 => UQVN_N97, A0 => A2, A1 => A1, A2 => A0, 
	A3 => UQVN_N146, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B126 : AND8
	PORT MAP (Z0 => UQVN_N95, A0 => A3, A1 => A1, A2 => A0, 
	A3 => UQVN_N145, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B127 : AND8
	PORT MAP (Z0 => UQVN_N96, A0 => A3, A1 => A2, A2 => A0, 
	A3 => UQVN_N144, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B128 : AND7
	PORT MAP (Z0 => UQVN_N106, A0 => A1, A1 => UQVN_N146, A2 => UQVN_N145, 
	A3 => UQVN_N144, A4 => UQVN_N116, A5 => UQVN_N148, A6 => UQVN_N115);
UQVB_B129 : AND8
	PORT MAP (Z0 => UQVN_N107, A0 => A3, A1 => A2, A2 => A1, 
	A3 => A0, A4 => UQVN_N143, A5 => UQVN_N116, A6 => UQVN_N148, 
	A7 => UQVN_N115);
UQVB_B130 : AND8
	PORT MAP (Z0 => UQVN_N123, A0 => UQVN_N142, A1 => UQVN_N139, A2 => B2, 
	A3 => B1, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B131 : AND8
	PORT MAP (Z0 => UQVN_N124, A0 => UQVN_N141, A1 => UQVN_N139, A2 => B3, 
	A3 => B1, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B132 : AND8
	PORT MAP (Z0 => UQVN_N125, A0 => UQVN_N140, A1 => UQVN_N139, A2 => B3, 
	A3 => B2, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B133 : AND8
	PORT MAP (Z0 => UQVN_N126, A0 => UQVN_N139, A1 => B3, A2 => B2, 
	A3 => B1, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B134 : AND7
	PORT MAP (Z0 => UQVN_N127, A0 => UQVN_N142, A1 => UQVN_N141, A2 => UQVN_N140, 
	A3 => B1, A4 => UQVN_N118, A5 => UQVN_N148, A6 => UQVN_N117);
UQVB_B135 : AND7
	PORT MAP (Z0 => UQVN_N128, A0 => UQVN_N142, A1 => UQVN_N140, A2 => B2, 
	A3 => B1, A4 => UQVN_N118, A5 => UQVN_N148, A6 => UQVN_N117);
UQVB_B136 : AND7
	PORT MAP (Z0 => UQVN_N129, A0 => UQVN_N141, A1 => UQVN_N140, A2 => B3, 
	A3 => B1, A4 => UQVN_N118, A5 => UQVN_N148, A6 => UQVN_N117);
UQVB_B137 : AND7
	PORT MAP (Z0 => UQVN_N130, A0 => UQVN_N140, A1 => B3, A2 => B2, 
	A3 => B1, A4 => UQVN_N118, A5 => UQVN_N148, A6 => UQVN_N117);
UQVB_B138 : OR7
	PORT MAP (Z0 => UQVN_N137, A0 => UQVN_N119, A1 => UQVN_N120, A2 => UQVN_N121, 
	A3 => UQVN_N122, A4 => UQVN_N123, A5 => UQVN_N124, A6 => UQVN_N125);
UQVB_B139 : OR5
	PORT MAP (Z0 => UQVN_N135, A0 => UQVN_N126, A1 => UQVN_N127, A2 => UQVN_N128, 
	A3 => UQVN_N129, A4 => UQVN_N130);
UQVB_B140 : AND3
	PORT MAP (Z0 => UQVN_N134, A0 => UQVN_N117, A1 => UQVN_N138, A2 => UQVN_N149);
UQVB_B141 : AND6
	PORT MAP (Z0 => UQVN_N133, A0 => UQVN_N142, A1 => UQVN_N141, A2 => B2, 
	A3 => UQVN_N118, A4 => UQVN_N148, A5 => UQVN_N117);
UQVB_B142 : AND6
	PORT MAP (Z0 => UQVN_N132, A0 => UQVN_N141, A1 => B3, A2 => B2, 
	A3 => UQVN_N118, A4 => UQVN_N148, A5 => UQVN_N117);
UQVB_B143 : AND5
	PORT MAP (Z0 => UQVN_N131, A0 => UQVN_N142, A1 => B3, A2 => UQVN_N118, 
	A3 => UQVN_N148, A4 => UQVN_N117);
UQVB_B144 : OR4
	PORT MAP (Z0 => UQVN_N136, A0 => UQVN_N134, A1 => UQVN_N133, A2 => UQVN_N132, 
	A3 => UQVN_N131);
UQVB_B145 : OR3
	PORT MAP (Z0 => LT, A0 => UQVN_N136, A1 => UQVN_N135, A2 => UQVN_N137);
UQVB_B146 : AND8
	PORT MAP (Z0 => UQVN_N119, A0 => UQVN_N142, A1 => UQVN_N141, A2 => UQVN_N140, 
	A3 => UQVN_N139, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B147 : INV
	PORT MAP (ZN0 => UQVN_N118, A0 => UQVN_N149);
UQVB_B148 : INV
	PORT MAP (ZN0 => UQVN_N138, A0 => UQVN_N148);
UQVB_B149 : AND8
	PORT MAP (Z0 => UQVN_N120, A0 => UQVN_N142, A1 => UQVN_N141, A2 => UQVN_N139, 
	A3 => B1, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B150 : INV
	PORT MAP (ZN0 => UQVN_N117, A0 => UQVN_N147);
UQVB_B151 : AND8
	PORT MAP (Z0 => UQVN_N121, A0 => UQVN_N142, A1 => UQVN_N140, A2 => UQVN_N139, 
	A3 => B2, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
UQVB_B152 : AND8
	PORT MAP (Z0 => UQVN_N122, A0 => UQVN_N141, A1 => UQVN_N140, A2 => UQVN_N139, 
	A3 => B3, A4 => B0, A5 => UQVN_N118, A6 => UQVN_N148, 
	A7 => UQVN_N117);
END lattice_arch;
-- VHDL netlist for MULT24
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MULT24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic
    );
END MULT24;


ARCHITECTURE lattice_arch OF MULT24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => A1);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => A1, A1 => B0, A2 => UQVN_N26);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => A0);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N25, A2 => B1);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N24, A2 => B1);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N23, A1 => A1, A2 => B0);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N4, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N25, A2 => B1, 
	A3 => UQVN_N27);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N23, A1 => A1, A2 => B1);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => UQVN_N26, A2 => B2);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => UQVN_N24, A2 => B2);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => A0, A1 => B0, A2 => B2);
UQVB_B14 : OR5
	PORT MAP (Z0 => Z2, A0 => UQVN_N7, A1 => UQVN_N6, A2 => UQVN_N5, 
	A3 => UQVN_N8, A4 => UQVN_N9);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => B2);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => B3);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => B0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => B1);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N23, A1 => A1, A2 => B3);
UQVB_B20 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => A1, A1 => UQVN_N26, A2 => UQVN_N27, 
	A3 => B3);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => A1, A1 => UQVN_N25, A2 => UQVN_N27, 
	A3 => B3);
UQVB_B22 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => A0, A1 => A1, A2 => B2, 
	A3 => B3);
UQVB_B23 : AND5
	PORT MAP (Z0 => UQVN_N18, A0 => A0, A1 => A1, A2 => B1, 
	A3 => B2, A4 => UQVN_N28);
UQVB_B24 : AND5
	PORT MAP (Z0 => UQVN_N21, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B1, A4 => B3);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N23, A1 => UQVN_N27, A2 => B3);
UQVB_B26 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => A0, A1 => A1, A2 => UQVN_N26, 
	A3 => B2);
UQVB_B27 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => A1, A1 => B0, A2 => B1, 
	A3 => UQVN_N27, A4 => B3);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N23, A1 => A1, A2 => B2, 
	A3 => UQVN_N28);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N23, A1 => UQVN_N24, A2 => B3);
UQVB_B30 : AND6
	PORT MAP (Z0 => UQVN_N15, A0 => A0, A1 => A1, A2 => B0, 
	A3 => B1, A4 => UQVN_N27, A5 => UQVN_N28);
UQVB_B31 : OR6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N15, A1 => UQVN_N14, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N12, A5 => UQVN_N13);
UQVB_B32 : LXOR2
	PORT MAP (Z0 => Z3, A0 => B3, A1 => UQVN_N16);
UQVB_B33 : OR4
	PORT MAP (Z0 => Z4, A0 => UQVN_N19, A1 => UQVN_N18, A2 => UQVN_N17, 
	A3 => UQVN_N20);
UQVB_B34 : OR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N22, A1 => UQVN_N21);
END lattice_arch;
-- VHDL netlist for PG1
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PG1 IS 
    PORT (
        GI1 : IN std_logic;
        PI1 : IN std_logic;
        PGI1 : IN std_logic;
        PGO1 : OUT std_logic
    );
END PG1;


ARCHITECTURE lattice_arch OF PG1 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => PI1, A1 => PGI1);
UQVB_B2 : OR2
	PORT MAP (Z0 => PGO1, A0 => GI1, A1 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for PG2
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PG2 IS 
    PORT (
        GI2 : IN std_logic;
        PI2 : IN std_logic;
        GI1 : IN std_logic;
        PI1 : IN std_logic;
        PGI1 : IN std_logic;
        PGO2 : OUT std_logic
    );
END PG2;


ARCHITECTURE lattice_arch OF PG2 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : OR3
	PORT MAP (Z0 => PGO2, A0 => GI2, A1 => UQVN_N1, A2 => UQVN_N2);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => PI2, A1 => PI1, A2 => PGI1);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => PI2, A1 => GI1);
END lattice_arch;
-- VHDL netlist for PG3
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PG3 IS 
    PORT (
        GI3 : IN std_logic;
        PI3 : IN std_logic;
        GI2 : IN std_logic;
        PI2 : IN std_logic;
        GI1 : IN std_logic;
        PI1 : IN std_logic;
        PGI1 : IN std_logic;
        PGO3 : OUT std_logic
    );
END PG3;


ARCHITECTURE lattice_arch OF PG3 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => PGO3, A0 => GI3, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => PI3, A1 => GI2);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => PI3, A1 => PI2, A2 => GI1);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => PI3, A1 => PI2, A2 => PI1, 
	A3 => PGI1);
END lattice_arch;
-- VHDL netlist for PG4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PG4 IS 
    PORT (
        GI4 : IN std_logic;
        PI4 : IN std_logic;
        GI3 : IN std_logic;
        PI3 : IN std_logic;
        GI2 : IN std_logic;
        PI2 : IN std_logic;
        GI1 : IN std_logic;
        PI1 : IN std_logic;
        PGI1 : IN std_logic;
        PGO4 : OUT std_logic
    );
END PG4;


ARCHITECTURE lattice_arch OF PG4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : OR5
	PORT MAP (Z0 => PGO4, A0 => GI4, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3, A4 => UQVN_N4);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => PI4, A1 => GI3);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => PI4, A1 => PI3, A2 => GI2);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => PI4, A1 => PI3, A2 => PI2, 
	A3 => GI1);
UQVB_B5 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => PI4, A1 => PI3, A2 => PI2, 
	A3 => PI1, A4 => PGI1);
END lattice_arch;

-- VHDL netlist for MULT44
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MULT44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic
    );
END MULT44;


ARCHITECTURE lattice_arch OF MULT44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 C5, G012, G345, H0,
	 H1, H2, H3, L0,
	 L1, L2, L3, L4,
	 L5, P345 : std_logic;


  COMPONENT MULT24
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic
    );
  END COMPONENT;

for all: MULT24 use  entity  lat_vhd.MULT24(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT F3ADD
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        CI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        G012 : OUT std_logic;
        P012 : OUT std_logic
    );
  END COMPONENT;

for all: F3ADD use  entity  lat_vhd.F3ADD(lattice_arch);


  COMPONENT PG1
    PORT (
        GI1 : IN std_logic;
        PI1 : IN std_logic;
        PGI1 : IN std_logic;
        PGO1 : OUT std_logic
    );
  END COMPONENT;

for all: PG1 use  entity  lat_vhd.PG1(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

    Z0 <= L0;
    Z1 <= L1;
UQVB_B1 : MULT24
	PORT MAP (Z0 => L0, Z1 => L1, Z2 => L2, Z3 => L3, 
	Z4 => L4, Z5 => L5, A0 => A0, A1 => A1, 
	B0 => B0, B1 => B1, B2 => B2, B3 => B3);
UQVB_B2 : MULT24
	PORT MAP (Z0 => H0, Z1 => H1, Z2 => H2, Z3 => H3, 
	Z4 => UQVN_N8, Z5 => UQVN_N2, A0 => A2, A1 => A3, 
	B0 => B0, B1 => B1, B2 => B2, B3 => B3);
UQVB_B3 : LXOR2
	PORT MAP (Z0 => Z2, A0 => L2, A1 => H0);
UQVB_B4 : F3ADD
	PORT MAP (Z0 => Z3, Z1 => Z4, Z2 => Z5, G012 => G345, 
	P012 => P345, A0 => L3, A1 => L4, A2 => L5, 
	B0 => H1, B1 => H2, B2 => H3, CI => G012);
UQVB_B5 : PG1
	PORT MAP (PGO1 => C5, GI1 => G345, PI1 => P345, PGI1 => G012);
UQVB_B6 : LXOR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N8, A1 => C5);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N1, A1 => UQVN_N8, A2 => C5);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => UQVN_N2);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => C5);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N7, A1 => UQVN_N2);
UQVB_B12 : OR3
	PORT MAP (Z0 => Z7, A0 => UQVN_N4, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B13 : AND2
	PORT MAP (Z0 => G012, A0 => H0, A1 => L2);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => UQVN_N8);
END lattice_arch;
-- VHDL netlist for MUX16
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX16 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX16;


ARCHITECTURE lattice_arch OF MUX16 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20 : std_logic;


  COMPONENT OR16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR16 use  entity  lat_vhd.OR16(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : OR16
	PORT MAP (Z0 => Z0, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N16, 
	A3 => UQVN_N15, A4 => UQVN_N14, A5 => UQVN_N8, A6 => UQVN_N7, 
	A7 => UQVN_N5, A8 => UQVN_N6, A9 => UQVN_N9, A10 => UQVN_N10, 
	A11 => UQVN_N11, A12 => UQVN_N12, A13 => UQVN_N13, A14 => UQVN_N17, 
	A15 => UQVN_N18);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S3);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S2);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S1);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N18, A0 => A15, A1 => S0, A2 => S1, 
	A3 => S2, A4 => S3);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N17, A0 => A14, A1 => UQVN_N4, A2 => S1, 
	A3 => S2, A4 => S3);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N13, A0 => A13, A1 => S0, A2 => UQVN_N3, 
	A3 => S2, A4 => S3);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => A12, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => S2, A4 => S3);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N11, A0 => A11, A1 => S0, A2 => S1, 
	A3 => UQVN_N2, A4 => S3);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => A10, A1 => UQVN_N4, A2 => S1, 
	A3 => UQVN_N2, A4 => S3);
UQVB_B12 : AND5
	PORT MAP (Z0 => UQVN_N9, A0 => A9, A1 => S0, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => S3);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => A8, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => S3);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => A7, A1 => S0, A2 => S1, 
	A3 => S2, A4 => UQVN_N1);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => A6, A1 => UQVN_N4, A2 => S1, 
	A3 => S2, A4 => UQVN_N1);
UQVB_B16 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => A5, A1 => S0, A2 => UQVN_N3, 
	A3 => S2, A4 => UQVN_N1);
UQVB_B17 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => A4, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => S2, A4 => UQVN_N1);
UQVB_B18 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => A3, A1 => S0, A2 => S1, 
	A3 => UQVN_N2, A4 => UQVN_N1);
UQVB_B19 : AND5
	PORT MAP (Z0 => UQVN_N16, A0 => A2, A1 => UQVN_N4, A2 => S1, 
	A3 => UQVN_N2, A4 => UQVN_N1);
UQVB_B20 : AND5
	PORT MAP (Z0 => UQVN_N19, A0 => A1, A1 => S0, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => UQVN_N1);
UQVB_B21 : AND5
	PORT MAP (Z0 => UQVN_N20, A0 => A0, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => UQVN_N1);
END lattice_arch;
-- VHDL netlist for MUX16E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX16E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX16E;


ARCHITECTURE lattice_arch OF MUX16E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20 : std_logic;


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT OR16
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR16 use  entity  lat_vhd.OR16(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND6
	PORT MAP (Z0 => UQVN_N18, A0 => A15, A1 => S0, A2 => S1, 
	A3 => S2, A4 => S3, A5 => EN);
UQVB_B2 : AND6
	PORT MAP (Z0 => UQVN_N17, A0 => A14, A1 => UQVN_N4, A2 => S1, 
	A3 => S2, A4 => S3, A5 => EN);
UQVB_B3 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => A13, A1 => S0, A2 => UQVN_N3, 
	A3 => S2, A4 => S3, A5 => EN);
UQVB_B4 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => A12, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => S2, A4 => S3, A5 => EN);
UQVB_B5 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => A11, A1 => S0, A2 => S1, 
	A3 => UQVN_N2, A4 => S3, A5 => EN);
UQVB_B6 : AND6
	PORT MAP (Z0 => UQVN_N10, A0 => A10, A1 => UQVN_N4, A2 => S1, 
	A3 => UQVN_N2, A4 => S3, A5 => EN);
UQVB_B7 : AND6
	PORT MAP (Z0 => UQVN_N9, A0 => A9, A1 => S0, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => S3, A5 => EN);
UQVB_B8 : AND6
	PORT MAP (Z0 => UQVN_N6, A0 => A8, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => S3, A5 => EN);
UQVB_B9 : AND6
	PORT MAP (Z0 => UQVN_N5, A0 => A7, A1 => S0, A2 => S1, 
	A3 => S2, A4 => UQVN_N1, A5 => EN);
UQVB_B10 : AND6
	PORT MAP (Z0 => UQVN_N7, A0 => A6, A1 => UQVN_N4, A2 => S1, 
	A3 => S2, A4 => UQVN_N1, A5 => EN);
UQVB_B11 : AND6
	PORT MAP (Z0 => UQVN_N8, A0 => A5, A1 => S0, A2 => UQVN_N3, 
	A3 => S2, A4 => UQVN_N1, A5 => EN);
UQVB_B12 : AND6
	PORT MAP (Z0 => UQVN_N14, A0 => A4, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => S2, A4 => UQVN_N1, A5 => EN);
UQVB_B13 : AND6
	PORT MAP (Z0 => UQVN_N15, A0 => A3, A1 => S0, A2 => S1, 
	A3 => UQVN_N2, A4 => UQVN_N1, A5 => EN);
UQVB_B14 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => A2, A1 => UQVN_N4, A2 => S1, 
	A3 => UQVN_N2, A4 => UQVN_N1, A5 => EN);
UQVB_B15 : AND6
	PORT MAP (Z0 => UQVN_N19, A0 => A1, A1 => S0, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => UQVN_N1, A5 => EN);
UQVB_B16 : AND6
	PORT MAP (Z0 => UQVN_N20, A0 => A0, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => UQVN_N2, A4 => UQVN_N1, A5 => EN);
UQVB_B17 : OR16
	PORT MAP (Z0 => Z0, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N16, 
	A3 => UQVN_N15, A4 => UQVN_N14, A5 => UQVN_N8, A6 => UQVN_N7, 
	A7 => UQVN_N5, A8 => UQVN_N6, A9 => UQVN_N9, A10 => UQVN_N10, 
	A11 => UQVN_N11, A12 => UQVN_N12, A13 => UQVN_N13, A14 => UQVN_N17, 
	A15 => UQVN_N18);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S3);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S2);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S1);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX2
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX2;


ARCHITECTURE lattice_arch OF MUX2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => A1, A1 => S0);
UQVB_B3 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX22
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX22 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END MUX22;


ARCHITECTURE lattice_arch OF MUX22 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => B1, A1 => S0);
UQVB_B3 : OR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => UQVN_N4);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX22E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX22E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END MUX22E;


ARCHITECTURE lattice_arch OF MUX22E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => UQVN_N1, A2 => EN);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => B1, A1 => S0, A2 => EN);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B5 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => UQVN_N4, A2 => EN);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0, A2 => EN);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX24
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        C0 : IN std_logic;
        C1 : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END MUX24;


ARCHITECTURE lattice_arch OF MUX24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N4);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => S0, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => C0, A1 => UQVN_N5, A2 => S1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => S0, A2 => S1);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S1);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N7, A1 => UQVN_N8, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N11, A2 => UQVN_N12);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => B1, A1 => S0, A2 => UQVN_N12);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => C1, A1 => UQVN_N11, A2 => S1);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D1, A1 => S0, A2 => S1);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => S1);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX24E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX24E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        C0 : IN std_logic;
        C1 : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic
    );
END MUX24E;


ARCHITECTURE lattice_arch OF MUX24E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N5);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => C0, A1 => UQVN_N4, A2 => S1, 
	A3 => EN);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N8, A1 => UQVN_N12, A2 => UQVN_N7, 
	A3 => UQVN_N11);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => S1);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => D1, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => C1, A1 => UQVN_N10, A2 => S1, 
	A3 => EN);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => B1, A1 => S0, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => A1, A1 => UQVN_N10, A2 => UQVN_N9, 
	A3 => EN);
END lattice_arch;
-- VHDL netlist for MUX2E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX2E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX2E;


ARCHITECTURE lattice_arch OF MUX2E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N1, A2 => EN);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => A1, A1 => S0, A2 => EN);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX4;


ARCHITECTURE lattice_arch OF MUX4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N4);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => S0, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => A2, A1 => UQVN_N5, A2 => S1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => A3, A1 => S0, A2 => S1);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S1);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX42
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX42 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END MUX42;


ARCHITECTURE lattice_arch OF MUX42 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => B1, A1 => S0);
UQVB_B3 : OR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => UQVN_N4);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => A3, A1 => UQVN_N7);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => B3, A1 => S0);
UQVB_B11 : OR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A2, A1 => UQVN_N10);
UQVB_B14 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => B2, A1 => S0);
UQVB_B15 : OR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX42E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX42E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END MUX42E;


ARCHITECTURE lattice_arch OF MUX42E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => A1, A1 => UQVN_N1, A2 => EN);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => B1, A1 => S0, A2 => EN);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B5 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A0, A1 => UQVN_N4, A2 => EN);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0, A2 => EN);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B9 : OR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A3, A1 => UQVN_N7, A2 => EN);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B3, A1 => S0, A2 => EN);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B13 : OR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => A2, A1 => UQVN_N10, A2 => EN);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => B2, A1 => S0, A2 => EN);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX44
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        C0 : IN std_logic;
        C1 : IN std_logic;
        C2 : IN std_logic;
        C3 : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END MUX44;


ARCHITECTURE lattice_arch OF MUX44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N4);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => S0, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => C0, A1 => UQVN_N5, A2 => S1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => S0, A2 => S1);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S1);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N7, A1 => UQVN_N8, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N11, A2 => UQVN_N12);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => B1, A1 => S0, A2 => UQVN_N12);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => C1, A1 => UQVN_N11, A2 => S1);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D1, A1 => S0, A2 => S1);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => S1);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => S0);
UQVB_B15 : OR4
	PORT MAP (Z0 => Z3, A0 => UQVN_N13, A1 => UQVN_N14, A2 => UQVN_N15, 
	A3 => UQVN_N16);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A3, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => B3, A1 => S0, A2 => UQVN_N18);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => C3, A1 => UQVN_N17, A2 => S1);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => D3, A1 => S0, A2 => S1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => S1);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => S0);
UQVB_B22 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N19, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N22);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => A2, A1 => UQVN_N23, A2 => UQVN_N24);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => B2, A1 => S0, A2 => UQVN_N24);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => C2, A1 => UQVN_N23, A2 => S1);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D2, A1 => S0, A2 => S1);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => S1);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX44A
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX44A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        C0 : IN std_logic;
        C1 : IN std_logic;
        C2 : IN std_logic;
        C3 : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END MUX44A;


ARCHITECTURE lattice_arch OF MUX44A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2, A2 => UQVN_N3, 
	A3 => UQVN_N4);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N5, A2 => UQVN_N6);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => S0, A2 => UQVN_N6);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => C0, A1 => UQVN_N5, A2 => S1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => D0, A1 => S0, A2 => S1);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S1);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S0);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N7, A1 => UQVN_N8, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N11, A2 => UQVN_N12);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => B1, A1 => S0, A2 => UQVN_N12);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => C1, A1 => UQVN_N11, A2 => S1);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => D1, A1 => S0, A2 => S1);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => S1);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => S0);
UQVB_B15 : OR4
	PORT MAP (Z0 => Z3, A0 => UQVN_N13, A1 => UQVN_N14, A2 => UQVN_N15, 
	A3 => UQVN_N16);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => A3, A1 => UQVN_N17, A2 => UQVN_N18);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => B3, A1 => S0, A2 => UQVN_N18);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => C3, A1 => UQVN_N17, A2 => S1);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => D3, A1 => S0, A2 => S1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => S1);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => S0);
UQVB_B22 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N19, A1 => UQVN_N20, A2 => UQVN_N21, 
	A3 => UQVN_N22);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => A2, A1 => UQVN_N23, A2 => UQVN_N24);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => B2, A1 => S0, A2 => UQVN_N24);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => C2, A1 => UQVN_N23, A2 => S1);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => D2, A1 => S0, A2 => S1);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => S1);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX44AE
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX44AE IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        C0 : IN std_logic;
        C1 : IN std_logic;
        C2 : IN std_logic;
        C3 : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END MUX44AE;


ARCHITECTURE lattice_arch OF MUX44AE IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N5);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => C0, A1 => UQVN_N4, A2 => S1, 
	A3 => EN);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N8, A1 => UQVN_N12, A2 => UQVN_N7, 
	A3 => UQVN_N11);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => S1);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => D1, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => C1, A1 => UQVN_N10, A2 => S1, 
	A3 => EN);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => B1, A1 => S0, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => A1, A1 => UQVN_N10, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B15 : OR4
	PORT MAP (Z0 => Z3, A0 => UQVN_N14, A1 => UQVN_N18, A2 => UQVN_N13, 
	A3 => UQVN_N17);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => S1);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => S0);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => D3, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => C3, A1 => UQVN_N16, A2 => S1, 
	A3 => EN);
UQVB_B20 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => B3, A1 => S0, A2 => UQVN_N15, 
	A3 => EN);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => A3, A1 => UQVN_N16, A2 => UQVN_N15, 
	A3 => EN);
UQVB_B22 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N20, A1 => UQVN_N24, A2 => UQVN_N19, 
	A3 => UQVN_N23);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => S1);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => S0);
UQVB_B25 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => D2, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B26 : AND4
	PORT MAP (Z0 => UQVN_N19, A0 => C2, A1 => UQVN_N22, A2 => S1, 
	A3 => EN);
UQVB_B27 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => B2, A1 => S0, A2 => UQVN_N21, 
	A3 => EN);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => A2, A1 => UQVN_N22, A2 => UQVN_N21, 
	A3 => EN);
END lattice_arch;
-- VHDL netlist for MUX44E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX44E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        C0 : IN std_logic;
        C1 : IN std_logic;
        C2 : IN std_logic;
        C3 : IN std_logic;
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END MUX44E;


ARCHITECTURE lattice_arch OF MUX44E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N5);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => D0, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => C0, A1 => UQVN_N4, A2 => S1, 
	A3 => EN);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => B0, A1 => S0, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B8 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N8, A1 => UQVN_N12, A2 => UQVN_N7, 
	A3 => UQVN_N11);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => S1);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => D1, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => C1, A1 => UQVN_N10, A2 => S1, 
	A3 => EN);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => B1, A1 => S0, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => A1, A1 => UQVN_N10, A2 => UQVN_N9, 
	A3 => EN);
UQVB_B15 : OR4
	PORT MAP (Z0 => Z3, A0 => UQVN_N14, A1 => UQVN_N18, A2 => UQVN_N13, 
	A3 => UQVN_N17);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => S1);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => S0);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => D3, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => C3, A1 => UQVN_N16, A2 => S1, 
	A3 => EN);
UQVB_B20 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => B3, A1 => S0, A2 => UQVN_N15, 
	A3 => EN);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => A3, A1 => UQVN_N16, A2 => UQVN_N15, 
	A3 => EN);
UQVB_B22 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N20, A1 => UQVN_N24, A2 => UQVN_N19, 
	A3 => UQVN_N23);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => S1);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => S0);
UQVB_B25 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => D2, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B26 : AND4
	PORT MAP (Z0 => UQVN_N19, A0 => C2, A1 => UQVN_N22, A2 => S1, 
	A3 => EN);
UQVB_B27 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => B2, A1 => S0, A2 => UQVN_N21, 
	A3 => EN);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => A2, A1 => UQVN_N22, A2 => UQVN_N21, 
	A3 => EN);
END lattice_arch;
-- VHDL netlist for MUX4E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX4E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX4E;


ARCHITECTURE lattice_arch OF MUX4E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N6, A2 => UQVN_N1, 
	A3 => UQVN_N5);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => A3, A1 => S0, A2 => S1, 
	A3 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N1, A0 => A2, A1 => UQVN_N4, A2 => S1, 
	A3 => EN);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => A1, A1 => S0, A2 => UQVN_N3, 
	A3 => EN);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => EN);
END lattice_arch;
-- VHDL netlist for MUX8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX8;


ARCHITECTURE lattice_arch OF MUX8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11 : std_logic;


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR8
	PORT MAP (Z0 => Z0, A0 => UQVN_N4, A1 => UQVN_N5, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8, A5 => UQVN_N11, A6 => UQVN_N10, 
	A7 => UQVN_N9);
UQVB_B2 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => A0, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B3 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => A1, A1 => S0, A2 => UQVN_N2, 
	A3 => UQVN_N3);
UQVB_B4 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => A2, A1 => UQVN_N1, A2 => S1, 
	A3 => UQVN_N3);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N7, A0 => A3, A1 => S0, A2 => S1, 
	A3 => UQVN_N3);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => A4, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => S2);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => A7, A1 => S0, A2 => S1, 
	A3 => S2);
UQVB_B8 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => A6, A1 => UQVN_N1, A2 => S1, 
	A3 => S2);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B10 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A5, A1 => S0, A2 => UQVN_N2, 
	A3 => S2);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S2);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
END lattice_arch;
-- VHDL netlist for MUX82
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX82 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic
    );
END MUX82;


ARCHITECTURE lattice_arch OF MUX82 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N1);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => B0, A1 => S0);
UQVB_B3 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => A1, A1 => UQVN_N4);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => B1, A1 => S0);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => A2, A1 => UQVN_N7);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => B2, A1 => S0);
UQVB_B11 : OR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => A3, A1 => UQVN_N10);
UQVB_B14 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => B3, A1 => S0);
UQVB_B15 : OR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => A4, A1 => UQVN_N13);
UQVB_B18 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => B4, A1 => S0);
UQVB_B19 : OR2
	PORT MAP (Z0 => Z4, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => S0);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => A5, A1 => UQVN_N16);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => B5, A1 => S0);
UQVB_B23 : OR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N17, A1 => UQVN_N18);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => S0);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => A6, A1 => UQVN_N19);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => B6, A1 => S0);
UQVB_B27 : OR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N20, A1 => UQVN_N21);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => S0);
UQVB_B29 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => A7, A1 => UQVN_N22);
UQVB_B30 : AND2
	PORT MAP (Z0 => UQVN_N24, A0 => B7, A1 => S0);
UQVB_B31 : OR2
	PORT MAP (Z0 => Z7, A0 => UQVN_N23, A1 => UQVN_N24);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX82E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX82E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic
    );
END MUX82E;


ARCHITECTURE lattice_arch OF MUX82E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => UQVN_N1, A2 => EN);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => B0, A1 => S0, A2 => EN);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B5 : OR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N5, A1 => UQVN_N6);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => A1, A1 => UQVN_N4, A2 => EN);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => B1, A1 => S0, A2 => EN);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => S0);
UQVB_B9 : OR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N8, A1 => UQVN_N9);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A2, A1 => UQVN_N7, A2 => EN);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B2, A1 => S0, A2 => EN);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S0);
UQVB_B13 : OR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => A3, A1 => UQVN_N10, A2 => EN);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => B3, A1 => S0, A2 => EN);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => S0);
UQVB_B17 : OR2
	PORT MAP (Z0 => Z4, A0 => UQVN_N14, A1 => UQVN_N15);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => A4, A1 => UQVN_N13, A2 => EN);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => B4, A1 => S0, A2 => EN);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => S0);
UQVB_B21 : OR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N17, A1 => UQVN_N18);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => A5, A1 => UQVN_N16, A2 => EN);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => B5, A1 => S0, A2 => EN);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => S0);
UQVB_B25 : OR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N20, A1 => UQVN_N21);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => A6, A1 => UQVN_N19, A2 => EN);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N21, A0 => B6, A1 => S0, A2 => EN);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => S0);
UQVB_B29 : OR2
	PORT MAP (Z0 => Z7, A0 => UQVN_N23, A1 => UQVN_N24);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => A7, A1 => UQVN_N22, A2 => EN);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => B7, A1 => S0, A2 => EN);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => S0);
END lattice_arch;
-- VHDL netlist for MUX8E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY MUX8E IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        EN : IN std_logic;
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        Z0 : OUT std_logic
    );
END MUX8E;


ARCHITECTURE lattice_arch OF MUX8E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11 : std_logic;


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : OR8
	PORT MAP (Z0 => Z0, A0 => UQVN_N4, A1 => UQVN_N5, A2 => UQVN_N6, 
	A3 => UQVN_N7, A4 => UQVN_N8, A5 => UQVN_N11, A6 => UQVN_N10, 
	A7 => UQVN_N9);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S0);
UQVB_B3 : AND5
	PORT MAP (Z0 => UQVN_N9, A0 => A7, A1 => S0, A2 => S1, 
	A3 => S2, A4 => EN);
UQVB_B4 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => A6, A1 => UQVN_N1, A2 => S1, 
	A3 => S2, A4 => EN);
UQVB_B5 : AND5
	PORT MAP (Z0 => UQVN_N11, A0 => A5, A1 => S0, A2 => UQVN_N2, 
	A3 => S2, A4 => EN);
UQVB_B6 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => A4, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => S2, A4 => EN);
UQVB_B7 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => A3, A1 => S0, A2 => S1, 
	A3 => UQVN_N3, A4 => EN);
UQVB_B8 : AND5
	PORT MAP (Z0 => UQVN_N6, A0 => A2, A1 => UQVN_N1, A2 => S1, 
	A3 => UQVN_N3, A4 => EN);
UQVB_B9 : AND5
	PORT MAP (Z0 => UQVN_N5, A0 => A1, A1 => S0, A2 => UQVN_N2, 
	A3 => UQVN_N3, A4 => EN);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => S2);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => A0, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => UQVN_N3, A4 => EN);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
END lattice_arch;
-- VHDL netlist for OB11
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OB11 IS 
    PORT (
        A0 : IN std_logic;
        XO0 : OUT std_logic
    );
END OB11;


ARCHITECTURE lattice_arch OF OB11 IS

  COMPONENT XOUTPUT
    PORT (
        A0 : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XOUTPUT use  entity  lat_vhd.XOUTPUT(lattice_arch);


BEGIN

UQVB_B1 : XOUTPUT
	PORT MAP (XO0 => XO0, A0 => A0);
END lattice_arch;
-- VHDL netlist for OB21
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OB21 IS 
    PORT (
        A0 : IN std_logic;
        XO0 : OUT std_logic
    );
END OB21;


ARCHITECTURE lattice_arch OF OB21 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XOUTPUT
    PORT (
        A0 : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XOUTPUT use  entity  lat_vhd.XOUTPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XOUTPUT
	PORT MAP (XO0 => XO0, A0 => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
END lattice_arch;
-- VHDL netlist for OB24
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OB24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic
    );
END OB24;


ARCHITECTURE lattice_arch OF OB24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XOUTPUT
    PORT (
        A0 : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XOUTPUT use  entity  lat_vhd.XOUTPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XOUTPUT
	PORT MAP (XO0 => XO3, A0 => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XOUTPUT
	PORT MAP (XO0 => XO2, A0 => UQVN_N2);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A2);
UQVB_B5 : XOUTPUT
	PORT MAP (XO0 => XO1, A0 => UQVN_N3);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A1);
UQVB_B7 : XOUTPUT
	PORT MAP (XO0 => XO0, A0 => UQVN_N4);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
END lattice_arch;
-- VHDL netlist for OB28
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OB28 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic;
        XO4 : OUT std_logic;
        XO5 : OUT std_logic;
        XO6 : OUT std_logic;
        XO7 : OUT std_logic
    );
END OB28;


ARCHITECTURE lattice_arch OF OB28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XOUTPUT
    PORT (
        A0 : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XOUTPUT use  entity  lat_vhd.XOUTPUT(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XOUTPUT
	PORT MAP (XO0 => XO6, A0 => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A6);
UQVB_B3 : XOUTPUT
	PORT MAP (XO0 => XO4, A0 => UQVN_N2);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A4);
UQVB_B5 : XOUTPUT
	PORT MAP (XO0 => XO2, A0 => UQVN_N3);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A2);
UQVB_B7 : XOUTPUT
	PORT MAP (XO0 => XO0, A0 => UQVN_N4);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
UQVB_B9 : XOUTPUT
	PORT MAP (XO0 => XO1, A0 => UQVN_N5);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A1);
UQVB_B11 : XOUTPUT
	PORT MAP (XO0 => XO3, A0 => UQVN_N6);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A3);
UQVB_B13 : XOUTPUT
	PORT MAP (XO0 => XO5, A0 => UQVN_N7);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A5);
UQVB_B15 : XOUTPUT
	PORT MAP (XO0 => XO7, A0 => UQVN_N8);
UQVB_B16 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A7);
END lattice_arch;
-- VHDL netlist for OT11
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT11 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
END OT11;


ARCHITECTURE lattice_arch OF OT11 IS

  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for OT14
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT14 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic
    );
END OT14;


ARCHITECTURE lattice_arch OF OT14 IS

  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => A3, OE => OE);
UQVB_B2 : XTRI1
	PORT MAP (XO0 => XO2, A0 => A2, OE => OE);
UQVB_B3 : XTRI1
	PORT MAP (XO0 => XO1, A0 => A1, OE => OE);
UQVB_B4 : XTRI1
	PORT MAP (XO0 => XO0, A0 => A0, OE => OE);
END lattice_arch;
-- VHDL netlist for OT18
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT18 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic;
        XO4 : OUT std_logic;
        XO5 : OUT std_logic;
        XO6 : OUT std_logic;
        XO7 : OUT std_logic
    );
END OT18;


ARCHITECTURE lattice_arch OF OT18 IS

  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => A3, OE => OE);
UQVB_B2 : XTRI1
	PORT MAP (XO0 => XO2, A0 => A2, OE => OE);
UQVB_B3 : XTRI1
	PORT MAP (XO0 => XO1, A0 => A1, OE => OE);
UQVB_B4 : XTRI1
	PORT MAP (XO0 => XO0, A0 => A0, OE => OE);
UQVB_B5 : XTRI1
	PORT MAP (XO0 => XO4, A0 => A4, OE => OE);
UQVB_B6 : XTRI1
	PORT MAP (XO0 => XO5, A0 => A5, OE => OE);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO6, A0 => A6, OE => OE);
UQVB_B8 : XTRI1
	PORT MAP (XO0 => XO7, A0 => A7, OE => OE);
END lattice_arch;
-- VHDL netlist for OT21
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT21 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
END OT21;


ARCHITECTURE lattice_arch OF OT21 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO0, A0 => UQVN_N1, OE => OE);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
END lattice_arch;
-- VHDL netlist for OT24
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT24 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic
    );
END OT24;


ARCHITECTURE lattice_arch OF OT24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => UQVN_N1, OE => OE);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XTRI1
	PORT MAP (XO0 => XO2, A0 => UQVN_N2, OE => OE);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A2);
UQVB_B5 : XTRI1
	PORT MAP (XO0 => XO1, A0 => UQVN_N3, OE => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A1);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO0, A0 => UQVN_N4, OE => OE);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
END lattice_arch;
-- VHDL netlist for OT28
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT28 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic;
        XO4 : OUT std_logic;
        XO5 : OUT std_logic;
        XO6 : OUT std_logic;
        XO7 : OUT std_logic
    );
END OT28;


ARCHITECTURE lattice_arch OF OT28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => UQVN_N1, OE => OE);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => A3);
UQVB_B3 : XTRI1
	PORT MAP (XO0 => XO2, A0 => UQVN_N2, OE => OE);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A2);
UQVB_B5 : XTRI1
	PORT MAP (XO0 => XO1, A0 => UQVN_N3, OE => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => A1);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO0, A0 => UQVN_N4, OE => OE);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
UQVB_B9 : XTRI1
	PORT MAP (XO0 => XO4, A0 => UQVN_N5, OE => OE);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => A4);
UQVB_B11 : XTRI1
	PORT MAP (XO0 => XO5, A0 => UQVN_N6, OE => OE);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A5);
UQVB_B13 : XTRI1
	PORT MAP (XO0 => XO6, A0 => UQVN_N7, OE => OE);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => A6);
UQVB_B15 : XTRI1
	PORT MAP (XO0 => XO7, A0 => UQVN_N8, OE => OE);
UQVB_B16 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A7);
END lattice_arch;
-- VHDL netlist for OT31
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT31 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
END OT31;


ARCHITECTURE lattice_arch OF OT31 IS
SIGNAL  UQVN_N1 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO0, A0 => A0, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
END lattice_arch;
-- VHDL netlist for OT34
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT34 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic
    );
END OT34;


ARCHITECTURE lattice_arch OF OT34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => A3, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XTRI1
	PORT MAP (XO0 => XO2, A0 => A2, OE => UQVN_N2);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B5 : XTRI1
	PORT MAP (XO0 => XO1, A0 => A1, OE => UQVN_N3);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO0, A0 => A0, OE => UQVN_N4);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
END lattice_arch;
-- VHDL netlist for OT38
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT38 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic;
        XO4 : OUT std_logic;
        XO5 : OUT std_logic;
        XO6 : OUT std_logic;
        XO7 : OUT std_logic
    );
END OT38;


ARCHITECTURE lattice_arch OF OT38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => A3, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XTRI1
	PORT MAP (XO0 => XO2, A0 => A2, OE => UQVN_N2);
UQVB_B4 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => OE);
UQVB_B5 : XTRI1
	PORT MAP (XO0 => XO1, A0 => A1, OE => UQVN_N3);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO0, A0 => A0, OE => UQVN_N4);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => OE);
UQVB_B9 : XTRI1
	PORT MAP (XO0 => XO4, A0 => A4, OE => UQVN_N5);
UQVB_B10 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => OE);
UQVB_B11 : XTRI1
	PORT MAP (XO0 => XO5, A0 => A5, OE => UQVN_N6);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => OE);
UQVB_B13 : XTRI1
	PORT MAP (XO0 => XO6, A0 => A6, OE => UQVN_N7);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => OE);
UQVB_B15 : XTRI1
	PORT MAP (XO0 => XO7, A0 => A7, OE => UQVN_N8);
UQVB_B16 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => OE);
END lattice_arch;
-- VHDL netlist for OT41
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT41 IS 
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
END OT41;


ARCHITECTURE lattice_arch OF OT41 IS
SIGNAL  UQVN_N1, UQVN_N2 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO0, A0 => UQVN_N2, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A0);
END lattice_arch;
-- VHDL netlist for OT44
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT44 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic
    );
END OT44;


ARCHITECTURE lattice_arch OF OT44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => UQVN_N2, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A3);
UQVB_B4 : XTRI1
	PORT MAP (XO0 => XO2, A0 => UQVN_N4, OE => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO1, A0 => UQVN_N6, OE => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => OE);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A1);
UQVB_B10 : XTRI1
	PORT MAP (XO0 => XO0, A0 => UQVN_N8, OE => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => OE);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A0);
END lattice_arch;
-- VHDL netlist for OT48
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY OT48 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic;
        XO1 : OUT std_logic;
        XO2 : OUT std_logic;
        XO3 : OUT std_logic;
        XO4 : OUT std_logic;
        XO5 : OUT std_logic;
        XO6 : OUT std_logic;
        XO7 : OUT std_logic
    );
END OT48;


ARCHITECTURE lattice_arch OF OT48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT XTRI1
    PORT (
        A0 : IN std_logic;
        OE : IN std_logic;
        XO0 : OUT std_logic
    );
  END COMPONENT;

for all: XTRI1 use  entity  lat_vhd.XTRI1(lattice_arch);


  COMPONENT XINV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: XINV use  entity  lat_vhd.XINV(lattice_arch);


BEGIN

UQVB_B1 : XTRI1
	PORT MAP (XO0 => XO3, A0 => UQVN_N2, OE => UQVN_N1);
UQVB_B2 : XINV
	PORT MAP (ZN0 => UQVN_N1, A0 => OE);
UQVB_B3 : XINV
	PORT MAP (ZN0 => UQVN_N2, A0 => A3);
UQVB_B4 : XTRI1
	PORT MAP (XO0 => XO2, A0 => UQVN_N4, OE => UQVN_N3);
UQVB_B5 : XINV
	PORT MAP (ZN0 => UQVN_N3, A0 => OE);
UQVB_B6 : XINV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B7 : XTRI1
	PORT MAP (XO0 => XO1, A0 => UQVN_N6, OE => UQVN_N5);
UQVB_B8 : XINV
	PORT MAP (ZN0 => UQVN_N5, A0 => OE);
UQVB_B9 : XINV
	PORT MAP (ZN0 => UQVN_N6, A0 => A1);
UQVB_B10 : XTRI1
	PORT MAP (XO0 => XO0, A0 => UQVN_N8, OE => UQVN_N7);
UQVB_B11 : XINV
	PORT MAP (ZN0 => UQVN_N7, A0 => OE);
UQVB_B12 : XINV
	PORT MAP (ZN0 => UQVN_N8, A0 => A0);
UQVB_B13 : XTRI1
	PORT MAP (XO0 => XO4, A0 => UQVN_N10, OE => UQVN_N9);
UQVB_B14 : XINV
	PORT MAP (ZN0 => UQVN_N9, A0 => OE);
UQVB_B15 : XINV
	PORT MAP (ZN0 => UQVN_N10, A0 => A4);
UQVB_B16 : XTRI1
	PORT MAP (XO0 => XO5, A0 => UQVN_N12, OE => UQVN_N11);
UQVB_B17 : XINV
	PORT MAP (ZN0 => UQVN_N11, A0 => OE);
UQVB_B18 : XINV
	PORT MAP (ZN0 => UQVN_N12, A0 => A5);
UQVB_B19 : XTRI1
	PORT MAP (XO0 => XO6, A0 => UQVN_N14, OE => UQVN_N13);
UQVB_B20 : XINV
	PORT MAP (ZN0 => UQVN_N13, A0 => OE);
UQVB_B21 : XINV
	PORT MAP (ZN0 => UQVN_N14, A0 => A6);
UQVB_B22 : XTRI1
	PORT MAP (XO0 => XO7, A0 => UQVN_N16, OE => UQVN_N15);
UQVB_B23 : XINV
	PORT MAP (ZN0 => UQVN_N15, A0 => OE);
UQVB_B24 : XINV
	PORT MAP (ZN0 => UQVN_N16, A0 => A7);
END lattice_arch;
-- VHDL netlist for PREN10
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PREN10 IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        S4 : IN std_logic;
        S5 : IN std_logic;
        S6 : IN std_logic;
        S7 : IN std_logic;
        S8 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END PREN10;


ARCHITECTURE lattice_arch OF PREN10 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => Z3, A0 => S8, A1 => S7);
UQVB_B2 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N1, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => UQVN_N2);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => S8);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S7);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N5, A1 => UQVN_N6, A2 => S3);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N6, A2 => S4);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N5, A1 => UQVN_N6, A2 => S5);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N5, A1 => UQVN_N6, A2 => S6);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N5, A1 => UQVN_N6, A2 => S5);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N5, A1 => UQVN_N6, A2 => S6);
UQVB_B11 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N9, A1 => UQVN_N8, A2 => UQVN_N10, 
	A3 => UQVN_N11);
UQVB_B12 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N5, A1 => UQVN_N6, A2 => UQVN_N12, 
	A3 => UQVN_N13, A4 => S2);
UQVB_B13 : AND5
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N5, A1 => UQVN_N6, A2 => UQVN_N12, 
	A3 => UQVN_N13, A4 => S1);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => S4);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => S3);
UQVB_B16 : OR5
	PORT MAP (Z0 => Z0, A0 => S8, A1 => UQVN_N14, A2 => UQVN_N15, 
	A3 => UQVN_N16, A4 => UQVN_N17);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N6, A1 => S6);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S4);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N6, A1 => UQVN_N7, A2 => UQVN_N13, 
	A3 => S2);
UQVB_B20 : AND5
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N6, A1 => UQVN_N7, A2 => UQVN_N13, 
	A3 => UQVN_N18, A4 => S0);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S5);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => S1);
END lattice_arch;
-- VHDL netlist for PREN10E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PREN10E IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        S4 : IN std_logic;
        S5 : IN std_logic;
        S6 : IN std_logic;
        S7 : IN std_logic;
        S8 : IN std_logic;
        EN : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END PREN10E;


ARCHITECTURE lattice_arch OF PREN10E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21 : std_logic;


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : OR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N20, A1 => UQVN_N21);
UQVB_B2 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N2, A1 => UQVN_N5, A2 => UQVN_N4, 
	A3 => UQVN_N3);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => S8);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => S7);
UQVB_B5 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N10, A1 => UQVN_N9, A2 => UQVN_N11, 
	A3 => UQVN_N12);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => S4);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => S3);
UQVB_B8 : OR5
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N15, A2 => UQVN_N16, 
	A3 => UQVN_N17, A4 => UQVN_N18);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => S5);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => S1);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => S8, A1 => EN);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => S7, A1 => EN);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S6, 
	A3 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S5, 
	A3 => EN);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S4, 
	A3 => EN);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S3, 
	A3 => EN);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S6, 
	A3 => EN);
UQVB_B18 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N6, A1 => UQVN_N7, A2 => S5, 
	A3 => EN);
UQVB_B19 : AND6
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N6, A1 => UQVN_N7, A2 => UQVN_N13, 
	A3 => UQVN_N14, A4 => S2, A5 => EN);
UQVB_B20 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N6, A1 => UQVN_N7, A2 => UQVN_N13, 
	A3 => UQVN_N14, A4 => S1, A5 => EN);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => S8, A1 => EN);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N7, A1 => S6, A2 => EN);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N7, A1 => UQVN_N8, A2 => S4, 
	A3 => EN);
UQVB_B24 : AND5
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N7, A1 => UQVN_N8, A2 => UQVN_N14, 
	A3 => S2, A4 => EN);
UQVB_B25 : AND6
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N7, A1 => UQVN_N8, A2 => UQVN_N14, 
	A3 => UQVN_N19, A4 => S0, A5 => EN);
END lattice_arch;
-- VHDL netlist for PREN16
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PREN16 IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        S4 : IN std_logic;
        S5 : IN std_logic;
        S6 : IN std_logic;
        S7 : IN std_logic;
        S8 : IN std_logic;
        S9 : IN std_logic;
        S10 : IN std_logic;
        S11 : IN std_logic;
        S12 : IN std_logic;
        S13 : IN std_logic;
        S14 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END PREN16;


ARCHITECTURE lattice_arch OF PREN16 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => S13);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => S12);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => S11);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => S10);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => S9);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => S8);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => S7);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => S5);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => S4);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => S3);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => S1);
UQVB_B12 : OR8
	PORT MAP (Z0 => Z3, A0 => S14, A1 => S13, A2 => S12, 
	A3 => S11, A4 => S10, A5 => S9, A6 => S8, 
	A7 => S7);
UQVB_B13 : OR8
	PORT MAP (Z0 => Z2, A0 => S14, A1 => S13, A2 => S12, 
	A3 => S11, A4 => UQVN_N1, A5 => UQVN_N2, A6 => UQVN_N3, 
	A7 => UQVN_N4);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N19, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => S6);
UQVB_B15 : AND5
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N19, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => S5);
UQVB_B16 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N19, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => S4);
UQVB_B17 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N19, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => S3);
UQVB_B18 : AND7
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N22, A1 => UQVN_N20, A2 => UQVN_N28, 
	A3 => UQVN_N26, A4 => UQVN_N25, A5 => UQVN_N23, A6 => S2);
UQVB_B19 : AND6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N22, A1 => UQVN_N20, A2 => UQVN_N28, 
	A3 => UQVN_N26, A4 => UQVN_N25, A5 => S4);
UQVB_B20 : AND5
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N22, A1 => UQVN_N20, A2 => UQVN_N28, 
	A3 => UQVN_N26, A4 => S6);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N22, A1 => UQVN_N20, A2 => UQVN_N28, 
	A3 => S8);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N22, A1 => UQVN_N20, A2 => S10);
UQVB_B23 : AND7
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N21, A1 => UQVN_N20, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => UQVN_N24, A5 => UQVN_N23, A6 => S1);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N21, A1 => UQVN_N20, A2 => S9);
UQVB_B25 : AND5
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N21, A1 => UQVN_N20, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => S6);
UQVB_B26 : AND7
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N21, A1 => UQVN_N20, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => UQVN_N24, A5 => UQVN_N23, A6 => S2);
UQVB_B27 : AND5
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N21, A1 => UQVN_N20, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => S5);
UQVB_B28 : OR8
	PORT MAP (Z0 => Z1, A0 => S14, A1 => S13, A2 => UQVN_N10, 
	A3 => UQVN_N9, A4 => UQVN_N8, A5 => UQVN_N7, A6 => UQVN_N6, 
	A7 => UQVN_N5);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N21, A1 => UQVN_N20, A2 => S10);
UQVB_B30 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N22, A1 => S12);
UQVB_B31 : OR8
	PORT MAP (Z0 => Z0, A0 => S14, A1 => UQVN_N11, A2 => UQVN_N17, 
	A3 => UQVN_N16, A4 => UQVN_N15, A5 => UQVN_N14, A6 => UQVN_N13, 
	A7 => UQVN_N12);
UQVB_B32 : AND8
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N22, A1 => UQVN_N20, A2 => UQVN_N28, 
	A3 => UQVN_N26, A4 => UQVN_N25, A5 => UQVN_N23, A6 => UQVN_N18, 
	A7 => S0);
END lattice_arch;
-- VHDL netlist for PREN16E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PREN16E IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        S4 : IN std_logic;
        S5 : IN std_logic;
        S6 : IN std_logic;
        S7 : IN std_logic;
        S8 : IN std_logic;
        S9 : IN std_logic;
        S10 : IN std_logic;
        S11 : IN std_logic;
        S12 : IN std_logic;
        S13 : IN std_logic;
        S14 : IN std_logic;
        EN : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic
    );
END PREN16E;


ARCHITECTURE lattice_arch OF PREN16E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => S13);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => S12);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => S11);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => S10);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => S9);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => S8);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => S7);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => S5);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => S4);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => S3);
UQVB_B11 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => S1);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => S14, A1 => EN);
UQVB_B13 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => S13, A1 => EN);
UQVB_B14 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => S12, A1 => EN);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => S11, A1 => EN);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => S10, A1 => EN);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => S9, A1 => EN);
UQVB_B18 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => S8, A1 => EN);
UQVB_B19 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => S7, A1 => EN);
UQVB_B20 : OR8
	PORT MAP (Z0 => Z3, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N2, A4 => UQVN_N1, A5 => UQVN_N3, A6 => UQVN_N4, 
	A7 => UQVN_N5);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N9, A0 => S11, A1 => EN);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N10, A0 => S12, A1 => EN);
UQVB_B23 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => S13, A1 => EN);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => S14, A1 => EN);
UQVB_B25 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N34, A1 => UQVN_N43, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => S6, A5 => EN);
UQVB_B26 : AND6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N34, A1 => UQVN_N43, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => S5, A5 => EN);
UQVB_B27 : AND6
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N34, A1 => UQVN_N43, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => S4, A5 => EN);
UQVB_B28 : AND6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N34, A1 => UQVN_N43, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => S3, A5 => EN);
UQVB_B29 : OR8
	PORT MAP (Z0 => Z2, A0 => UQVN_N12, A1 => UQVN_N11, A2 => UQVN_N10, 
	A3 => UQVN_N9, A4 => UQVN_N13, A5 => UQVN_N14, A6 => UQVN_N15, 
	A7 => UQVN_N16);
UQVB_B30 : AND9
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N37, A1 => UQVN_N35, A2 => UQVN_N43, 
	A3 => UQVN_N41, A4 => UQVN_N40, A5 => UQVN_N38, A6 => UQVN_N33, 
	A7 => S0, A8 => EN);
UQVB_B31 : AND8
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N37, A1 => UQVN_N35, A2 => UQVN_N43, 
	A3 => UQVN_N41, A4 => UQVN_N40, A5 => UQVN_N38, A6 => S2, 
	A7 => EN);
UQVB_B32 : AND7
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N37, A1 => UQVN_N35, A2 => UQVN_N43, 
	A3 => UQVN_N41, A4 => UQVN_N40, A5 => S4, A6 => EN);
UQVB_B33 : AND6
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N37, A1 => UQVN_N35, A2 => UQVN_N43, 
	A3 => UQVN_N41, A4 => S6, A5 => EN);
UQVB_B34 : AND5
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N37, A1 => UQVN_N35, A2 => UQVN_N43, 
	A3 => S8, A4 => EN);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N37, A1 => UQVN_N35, A2 => S10, 
	A3 => EN);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N37, A1 => S12, A2 => EN);
UQVB_B37 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => S14, A1 => EN);
UQVB_B38 : OR8
	PORT MAP (Z0 => Z0, A0 => UQVN_N17, A1 => UQVN_N24, A2 => UQVN_N18, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => UQVN_N21, A6 => UQVN_N22, 
	A7 => UQVN_N23);
UQVB_B39 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => S14, A1 => EN);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => S13, A1 => EN);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N36, A1 => UQVN_N35, A2 => S10, 
	A3 => EN);
UQVB_B42 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N36, A1 => UQVN_N35, A2 => S9, 
	A3 => EN);
UQVB_B43 : AND6
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N36, A1 => UQVN_N35, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => S6, A5 => EN);
UQVB_B44 : AND6
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N36, A1 => UQVN_N35, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => S5, A5 => EN);
UQVB_B45 : AND8
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N36, A1 => UQVN_N35, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => UQVN_N39, A5 => UQVN_N38, A6 => S2, 
	A7 => EN);
UQVB_B46 : AND8
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N36, A1 => UQVN_N35, A2 => UQVN_N42, 
	A3 => UQVN_N41, A4 => UQVN_N39, A5 => UQVN_N38, A6 => S1, 
	A7 => EN);
UQVB_B47 : OR8
	PORT MAP (Z0 => Z1, A0 => UQVN_N28, A1 => UQVN_N27, A2 => UQVN_N26, 
	A3 => UQVN_N25, A4 => UQVN_N29, A5 => UQVN_N30, A6 => UQVN_N31, 
	A7 => UQVN_N32);
END lattice_arch;
-- VHDL netlist for PREN8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PREN8 IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        S4 : IN std_logic;
        S5 : IN std_logic;
        S6 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic
    );
END PREN8;


ARCHITECTURE lattice_arch OF PREN8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N9, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => S0);
UQVB_B2 : OR4
	PORT MAP (Z0 => Z0, A0 => S6, A1 => UQVN_N5, A2 => UQVN_N4, 
	A3 => UQVN_N3);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
UQVB_B4 : OR4
	PORT MAP (Z0 => Z1, A0 => S6, A1 => S5, A2 => UQVN_N6, 
	A3 => UQVN_N7);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N8, A1 => S1, A2 => UQVN_N1);
UQVB_B6 : OR4
	PORT MAP (Z0 => Z2, A0 => S6, A1 => S5, A2 => S4, 
	A3 => S3);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S3);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => S4);
UQVB_B9 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N8, A1 => S2, A2 => UQVN_N1);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N9, A1 => UQVN_N1, A2 => S2);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N9, A1 => S4);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => S5);
END lattice_arch;
-- VHDL netlist for PREN8E
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY PREN8E IS 
    PORT (
        S0 : IN std_logic;
        S1 : IN std_logic;
        S2 : IN std_logic;
        S3 : IN std_logic;
        S4 : IN std_logic;
        S5 : IN std_logic;
        S6 : IN std_logic;
        EN : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic
    );
END PREN8E;


ARCHITECTURE lattice_arch OF PREN8E IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16 : std_logic;


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : OR4
	PORT MAP (Z0 => Z0, A0 => UQVN_N11, A1 => UQVN_N12, A2 => UQVN_N13, 
	A3 => UQVN_N14);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => S1);
UQVB_B3 : OR4
	PORT MAP (Z0 => Z1, A0 => UQVN_N7, A1 => UQVN_N8, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B4 : OR4
	PORT MAP (Z0 => Z2, A0 => UQVN_N6, A1 => UQVN_N4, A2 => UQVN_N3, 
	A3 => UQVN_N5);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => S3);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => S4);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => S3);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => EN, A1 => S4);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => EN, A1 => S5);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => EN, A1 => S6);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => EN, A1 => S6);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => EN, A1 => S5);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N15, A1 => S2, A2 => UQVN_N1, 
	A3 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N15, A1 => S1, A2 => UQVN_N1, 
	A3 => EN);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => EN, A1 => S6);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N16, A1 => S4, A2 => EN);
UQVB_B17 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N16, A1 => UQVN_N1, A2 => S2, 
	A3 => EN);
UQVB_B18 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N16, A1 => UQVN_N1, A2 => UQVN_N2, 
	A3 => S0, A4 => EN);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => S5);
END lattice_arch;
-- VHDL netlist for SRR11
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR11 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END SRR11;


ARCHITECTURE lattice_arch OF SRR11 IS

  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => Q0, D0 => CAI, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for SRR14
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR14 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END SRR14;


ARCHITECTURE lattice_arch OF SRR14 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3 : std_logic;


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


BEGIN

UQVB_B1 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N1);
UQVB_B2 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N2);
UQVB_B3 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N3);
UQVB_B4 : FD21
	PORT MAP (Q0 => Q3, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B5 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B6 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B7 : FD21
	PORT MAP (Q0 => UQVN_N1, D0 => CAI, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for SRR18
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR18 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END SRR18;


ARCHITECTURE lattice_arch OF SRR18 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N2, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : FD21
	PORT MAP (Q0 => Q7, D0 => UQVN_N4, CLK => CLK, CD => CD);
UQVB_B3 : FD21
	PORT MAP (Q0 => UQVN_N4, D0 => UQVN_N3, CLK => CLK, CD => CD);
UQVB_B4 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N2, CLK => CLK, CD => CD);
UQVB_B5 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N6);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N7);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N1);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N2);
UQVB_B10 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N3);
UQVB_B11 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N4);
UQVB_B12 : FD21
	PORT MAP (Q0 => UQVN_N1, D0 => UQVN_N7, CLK => CLK, CD => CD);
UQVB_B13 : FD21
	PORT MAP (Q0 => UQVN_N7, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B14 : FD21
	PORT MAP (Q0 => UQVN_N6, D0 => UQVN_N5, CLK => CLK, CD => CD);
UQVB_B15 : FD21
	PORT MAP (Q0 => UQVN_N5, D0 => CAI, CLK => CLK, CD => CD);
END lattice_arch;
-- VHDL netlist for SRR21
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR21 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END SRR21;


ARCHITECTURE lattice_arch OF SRR21 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => CAI, A1 => EN);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B6 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N5);
END lattice_arch;
-- VHDL netlist for SRR24
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR24 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END SRR24;


ARCHITECTURE lattice_arch OF SRR24 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23 : std_logic;


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N21);
UQVB_B2 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N22);
UQVB_B3 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N23);
UQVB_B4 : FD21
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N23, A1 => EN);
UQVB_B6 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B8 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N5);
UQVB_B10 : FD21
	PORT MAP (Q0 => UQVN_N10, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N22, A1 => EN);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N9);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => EN);
UQVB_B14 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B15 : BUF
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N10);
UQVB_B16 : FD21
	PORT MAP (Q0 => UQVN_N15, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B17 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N21, A1 => EN);
UQVB_B18 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N15, A1 => UQVN_N14);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => EN);
UQVB_B20 : OR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N12, A1 => UQVN_N13);
UQVB_B21 : BUF
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N15);
UQVB_B22 : FD21
	PORT MAP (Q0 => UQVN_N20, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B23 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => CAI, A1 => EN);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => EN);
UQVB_B26 : OR2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N17, A1 => UQVN_N18);
UQVB_B27 : BUF
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N20);
END lattice_arch;
-- VHDL netlist for SRR28
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR28 IS 
    PORT (
        CAI : IN std_logic;
        CLK : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END SRR28;


ARCHITECTURE lattice_arch OF SRR28 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N5, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N41, A1 => EN);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N5, A1 => UQVN_N4);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B5 : OR2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B6 : BUF
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N5);
UQVB_B7 : FD21
	PORT MAP (Q0 => UQVN_N10, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N44, A1 => EN);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N10, A1 => UQVN_N9);
UQVB_B10 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => EN);
UQVB_B11 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N7, A1 => UQVN_N8);
UQVB_B12 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N10);
UQVB_B13 : FD21
	PORT MAP (Q0 => UQVN_N15, D0 => UQVN_N11, CLK => CLK, CD => CD);
UQVB_B14 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N43, A1 => EN);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N15, A1 => UQVN_N14);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => EN);
UQVB_B17 : OR2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N12, A1 => UQVN_N13);
UQVB_B18 : BUF
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N15);
UQVB_B19 : FD21
	PORT MAP (Q0 => UQVN_N20, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N42, A1 => EN);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N20, A1 => UQVN_N19);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => EN);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N17, A1 => UQVN_N18);
UQVB_B24 : BUF
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N20);
UQVB_B25 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N45);
UQVB_B26 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N46);
UQVB_B27 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N47);
UQVB_B28 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N41);
UQVB_B29 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N42);
UQVB_B30 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N43);
UQVB_B31 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N44);
UQVB_B32 : FD21
	PORT MAP (Q0 => UQVN_N25, D0 => UQVN_N21, CLK => CLK, CD => CD);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N47, A1 => EN);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N25, A1 => UQVN_N24);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => EN);
UQVB_B36 : OR2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N22, A1 => UQVN_N23);
UQVB_B37 : BUF
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N25);
UQVB_B38 : FD21
	PORT MAP (Q0 => UQVN_N30, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B39 : AND2
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N46, A1 => EN);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N30, A1 => UQVN_N29);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => EN);
UQVB_B42 : OR2
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N27, A1 => UQVN_N28);
UQVB_B43 : BUF
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N30);
UQVB_B44 : FD21
	PORT MAP (Q0 => UQVN_N35, D0 => UQVN_N31, CLK => CLK, CD => CD);
UQVB_B45 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N45, A1 => EN);
UQVB_B46 : AND2
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N35, A1 => UQVN_N34);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => EN);
UQVB_B48 : OR2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N32, A1 => UQVN_N33);
UQVB_B49 : BUF
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N35);
UQVB_B50 : FD21
	PORT MAP (Q0 => UQVN_N40, D0 => UQVN_N36, CLK => CLK, CD => CD);
UQVB_B51 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => CAI, A1 => EN);
UQVB_B52 : AND2
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N39);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => EN);
UQVB_B54 : OR2
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N37, A1 => UQVN_N38);
UQVB_B55 : BUF
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N40);
END lattice_arch;
-- VHDL netlist for SRR31
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR31 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
END SRR31;


ARCHITECTURE lattice_arch OF SRR31 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => UQVN_N2, A2 => CAI);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => LD, A1 => D0);
UQVB_B5 : OR4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N5, A2 => UQVN_N7, 
	A3 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LD);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for SRR34
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR34 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END SRR34;


ARCHITECTURE lattice_arch OF SRR34 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N31);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => LD, A1 => D3);
UQVB_B5 : OR4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N5, A2 => UQVN_N7, 
	A3 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LD);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B8 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N3);
UQVB_B9 : FD21
	PORT MAP (Q0 => UQVN_N10, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N10, A1 => UQVN_N9, A2 => UQVN_N11);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => EN, A1 => UQVN_N9, A2 => UQVN_N30);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => LD, A1 => D2);
UQVB_B13 : OR4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N13, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => PS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => LD);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => EN);
UQVB_B16 : BUF
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N10);
UQVB_B17 : FD21
	PORT MAP (Q0 => UQVN_N17, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N18);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => EN, A1 => UQVN_N16, A2 => UQVN_N29);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => LD, A1 => D1);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N21, 
	A3 => PS);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => LD);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => EN);
UQVB_B24 : BUF
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N17);
UQVB_B25 : FD21
	PORT MAP (Q0 => UQVN_N24, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N25);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => EN, A1 => UQVN_N23, A2 => CAI);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => LD, A1 => D0);
UQVB_B29 : OR4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N28, 
	A3 => PS);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => LD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => EN);
UQVB_B32 : BUF
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N24);
UQVB_B33 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N31);
UQVB_B34 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N30);
UQVB_B35 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N29);
END lattice_arch;
-- VHDL netlist for SRR38
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR38 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END SRR38;


ARCHITECTURE lattice_arch OF SRR38 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63 : std_logic;


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD21
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N1, CLK => CLK, CD => CD);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N63);
UQVB_B4 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => LD, A1 => D3);
UQVB_B5 : OR4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N5, A2 => UQVN_N7, 
	A3 => PS);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LD);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B8 : BUF
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N3);
UQVB_B9 : FD21
	PORT MAP (Q0 => UQVN_N10, D0 => UQVN_N8, CLK => CLK, CD => CD);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N10, A1 => UQVN_N9, A2 => UQVN_N11);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => EN, A1 => UQVN_N9, A2 => UQVN_N62);
UQVB_B12 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => LD, A1 => D2);
UQVB_B13 : OR4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N13, A1 => UQVN_N12, A2 => UQVN_N14, 
	A3 => PS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => LD);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => EN);
UQVB_B16 : BUF
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N10);
UQVB_B17 : FD21
	PORT MAP (Q0 => UQVN_N17, D0 => UQVN_N15, CLK => CLK, CD => CD);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N18);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => EN, A1 => UQVN_N16, A2 => UQVN_N61);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => LD, A1 => D1);
UQVB_B21 : OR4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N21, 
	A3 => PS);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => LD);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => EN);
UQVB_B24 : BUF
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N17);
UQVB_B25 : FD21
	PORT MAP (Q0 => UQVN_N24, D0 => UQVN_N22, CLK => CLK, CD => CD);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N25);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => EN, A1 => UQVN_N23, A2 => CAI);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => LD, A1 => D0);
UQVB_B29 : OR4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N28, 
	A3 => PS);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => LD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => EN);
UQVB_B32 : BUF
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N24);
UQVB_B33 : FD21
	PORT MAP (Q0 => UQVN_N31, D0 => UQVN_N29, CLK => CLK, CD => CD);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N31, A1 => UQVN_N30, A2 => UQVN_N32);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => EN, A1 => UQVN_N30, A2 => UQVN_N57);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N35, A0 => LD, A1 => D4);
UQVB_B37 : OR4
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N34, A1 => UQVN_N33, A2 => UQVN_N35, 
	A3 => PS);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => LD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => EN);
UQVB_B40 : BUF
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N31);
UQVB_B41 : FD21
	PORT MAP (Q0 => UQVN_N38, D0 => UQVN_N36, CLK => CLK, CD => CD);
UQVB_B42 : AND3
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N39);
UQVB_B43 : AND3
	PORT MAP (Z0 => UQVN_N40, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N60);
UQVB_B44 : AND2
	PORT MAP (Z0 => UQVN_N42, A0 => LD, A1 => D5);
UQVB_B45 : OR4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N41, A1 => UQVN_N40, A2 => UQVN_N42, 
	A3 => PS);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => LD);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => EN);
UQVB_B48 : BUF
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N38);
UQVB_B49 : FD21
	PORT MAP (Q0 => UQVN_N45, D0 => UQVN_N43, CLK => CLK, CD => CD);
UQVB_B50 : AND3
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N45, A1 => UQVN_N44, A2 => UQVN_N46);
UQVB_B51 : AND3
	PORT MAP (Z0 => UQVN_N47, A0 => EN, A1 => UQVN_N44, A2 => UQVN_N59);
UQVB_B52 : AND2
	PORT MAP (Z0 => UQVN_N49, A0 => LD, A1 => D6);
UQVB_B53 : OR4
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N48, A1 => UQVN_N47, A2 => UQVN_N49, 
	A3 => PS);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => LD);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => EN);
UQVB_B56 : BUF
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N45);
UQVB_B57 : FD21
	PORT MAP (Q0 => UQVN_N52, D0 => UQVN_N50, CLK => CLK, CD => CD);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N52, A1 => UQVN_N51, A2 => UQVN_N53);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N54, A0 => EN, A1 => UQVN_N51, A2 => UQVN_N58);
UQVB_B60 : AND2
	PORT MAP (Z0 => UQVN_N56, A0 => LD, A1 => D7);
UQVB_B61 : OR4
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N55, A1 => UQVN_N54, A2 => UQVN_N56, 
	A3 => PS);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => LD);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => EN);
UQVB_B64 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N52);
UQVB_B65 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N58);
UQVB_B66 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N59);
UQVB_B67 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N60);
UQVB_B68 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N61);
UQVB_B69 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N62);
UQVB_B70 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N63);
UQVB_B71 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N57);
END lattice_arch;
-- VHDL netlist for SRR41
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR41 IS 
    PORT (
        D0 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic
    );
END SRR41;


ARCHITECTURE lattice_arch OF SRR41 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N5, A2 => UQVN_N7, 
	A3 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N8);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N8, 
	A3 => CAI);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => LD, A1 => UQVN_N8, A2 => D0);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N3);
END lattice_arch;
-- VHDL netlist for SRR44
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR44 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END SRR44;


ARCHITECTURE lattice_arch OF SRR44 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N5, A2 => UQVN_N7, 
	A3 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N8);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N8, 
	A3 => UQVN_N35);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => LD, A1 => UQVN_N8, A2 => D3);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B9 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N3);
UQVB_B10 : FD11
	PORT MAP (Q0 => UQVN_N11, D0 => UQVN_N9, CLK => CLK);
UQVB_B11 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N15, 
	A3 => PS);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => LD);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N11, A1 => UQVN_N10, A2 => UQVN_N12, 
	A3 => UQVN_N16);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => EN, A1 => UQVN_N10, A2 => UQVN_N16, 
	A3 => UQVN_N34);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => LD, A1 => UQVN_N16, A2 => D2);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => CS);
UQVB_B18 : BUF
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N11);
UQVB_B19 : FD11
	PORT MAP (Q0 => UQVN_N19, D0 => UQVN_N17, CLK => CLK);
UQVB_B20 : OR4
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N22, A1 => UQVN_N21, A2 => UQVN_N23, 
	A3 => PS);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => LD);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => EN);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N19, A1 => UQVN_N18, A2 => UQVN_N20, 
	A3 => UQVN_N24);
UQVB_B24 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => EN, A1 => UQVN_N18, A2 => UQVN_N24, 
	A3 => UQVN_N33);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => LD, A1 => UQVN_N24, A2 => D1);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => CS);
UQVB_B27 : BUF
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N19);
UQVB_B28 : FD11
	PORT MAP (Q0 => UQVN_N27, D0 => UQVN_N25, CLK => CLK);
UQVB_B29 : OR4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N30, A1 => UQVN_N29, A2 => UQVN_N31, 
	A3 => PS);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => LD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => EN);
UQVB_B32 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N28, 
	A3 => UQVN_N32);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => EN, A1 => UQVN_N26, A2 => UQVN_N32, 
	A3 => CAI);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => LD, A1 => UQVN_N32, A2 => D0);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => CS);
UQVB_B36 : BUF
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N27);
UQVB_B37 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N33);
UQVB_B38 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N34);
UQVB_B39 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N35);
END lattice_arch;
-- VHDL netlist for SRR48
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRR48 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAI : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END SRR48;


ARCHITECTURE lattice_arch OF SRR48 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71 : std_logic;


  COMPONENT FD11
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD11 use  entity  lat_vhd.FD11(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


BEGIN

UQVB_B1 : FD11
	PORT MAP (Q0 => UQVN_N3, D0 => UQVN_N1, CLK => CLK);
UQVB_B2 : OR4
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N6, A1 => UQVN_N5, A2 => UQVN_N7, 
	A3 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => LD);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => EN);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N4, 
	A3 => UQVN_N8);
UQVB_B6 : AND4
	PORT MAP (Z0 => UQVN_N5, A0 => EN, A1 => UQVN_N2, A2 => UQVN_N8, 
	A3 => UQVN_N71);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => LD, A1 => UQVN_N8, A2 => D3);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => CS);
UQVB_B9 : BUF
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N3);
UQVB_B10 : FD11
	PORT MAP (Q0 => UQVN_N11, D0 => UQVN_N9, CLK => CLK);
UQVB_B11 : OR4
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N14, A1 => UQVN_N13, A2 => UQVN_N15, 
	A3 => PS);
UQVB_B12 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => LD);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => EN);
UQVB_B14 : AND4
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N11, A1 => UQVN_N10, A2 => UQVN_N12, 
	A3 => UQVN_N16);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => EN, A1 => UQVN_N10, A2 => UQVN_N16, 
	A3 => UQVN_N70);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => LD, A1 => UQVN_N16, A2 => D2);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N16, A0 => CS);
UQVB_B18 : BUF
	PORT MAP (Z0 => UQVN_N71, A0 => UQVN_N11);
UQVB_B19 : FD11
	PORT MAP (Q0 => UQVN_N19, D0 => UQVN_N17, CLK => CLK);
UQVB_B20 : OR4
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N22, A1 => UQVN_N21, A2 => UQVN_N23, 
	A3 => PS);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => LD);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => EN);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N19, A1 => UQVN_N18, A2 => UQVN_N20, 
	A3 => UQVN_N24);
UQVB_B24 : AND4
	PORT MAP (Z0 => UQVN_N21, A0 => EN, A1 => UQVN_N18, A2 => UQVN_N24, 
	A3 => UQVN_N69);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => LD, A1 => UQVN_N24, A2 => D1);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => CS);
UQVB_B27 : BUF
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N19);
UQVB_B28 : FD11
	PORT MAP (Q0 => UQVN_N27, D0 => UQVN_N25, CLK => CLK);
UQVB_B29 : OR4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N30, A1 => UQVN_N29, A2 => UQVN_N31, 
	A3 => PS);
UQVB_B30 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => LD);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => EN);
UQVB_B32 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N27, A1 => UQVN_N26, A2 => UQVN_N28, 
	A3 => UQVN_N32);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => EN, A1 => UQVN_N26, A2 => UQVN_N32, 
	A3 => CAI);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => LD, A1 => UQVN_N32, A2 => D0);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => CS);
UQVB_B36 : BUF
	PORT MAP (Z0 => UQVN_N69, A0 => UQVN_N27);
UQVB_B37 : FD11
	PORT MAP (Q0 => UQVN_N35, D0 => UQVN_N33, CLK => CLK);
UQVB_B38 : OR4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N39, 
	A3 => PS);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => LD);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => EN);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N35, A1 => UQVN_N34, A2 => UQVN_N36, 
	A3 => UQVN_N40);
UQVB_B42 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => EN, A1 => UQVN_N34, A2 => UQVN_N40, 
	A3 => UQVN_N65);
UQVB_B43 : AND3
	PORT MAP (Z0 => UQVN_N39, A0 => LD, A1 => UQVN_N40, A2 => D4);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CS);
UQVB_B45 : BUF
	PORT MAP (Z0 => UQVN_N68, A0 => UQVN_N35);
UQVB_B46 : FD11
	PORT MAP (Q0 => UQVN_N43, D0 => UQVN_N41, CLK => CLK);
UQVB_B47 : OR4
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N46, A1 => UQVN_N45, A2 => UQVN_N47, 
	A3 => PS);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => LD);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => EN);
UQVB_B50 : AND4
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N43, A1 => UQVN_N42, A2 => UQVN_N44, 
	A3 => UQVN_N48);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N45, A0 => EN, A1 => UQVN_N42, A2 => UQVN_N48, 
	A3 => UQVN_N68);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N47, A0 => LD, A1 => UQVN_N48, A2 => D5);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => CS);
UQVB_B54 : BUF
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N43);
UQVB_B55 : FD11
	PORT MAP (Q0 => UQVN_N51, D0 => UQVN_N49, CLK => CLK);
UQVB_B56 : OR4
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N54, A1 => UQVN_N53, A2 => UQVN_N55, 
	A3 => PS);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => LD);
UQVB_B58 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => EN);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N51, A1 => UQVN_N50, A2 => UQVN_N52, 
	A3 => UQVN_N56);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N53, A0 => EN, A1 => UQVN_N50, A2 => UQVN_N56, 
	A3 => UQVN_N67);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N55, A0 => LD, A1 => UQVN_N56, A2 => D6);
UQVB_B62 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => CS);
UQVB_B63 : BUF
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N51);
UQVB_B64 : FD11
	PORT MAP (Q0 => UQVN_N59, D0 => UQVN_N57, CLK => CLK);
UQVB_B65 : OR4
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N62, A1 => UQVN_N61, A2 => UQVN_N63, 
	A3 => PS);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N58, A0 => LD);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N60, A0 => EN);
UQVB_B68 : AND4
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N59, A1 => UQVN_N58, A2 => UQVN_N60, 
	A3 => UQVN_N64);
UQVB_B69 : AND4
	PORT MAP (Z0 => UQVN_N61, A0 => EN, A1 => UQVN_N58, A2 => UQVN_N64, 
	A3 => UQVN_N66);
UQVB_B70 : AND3
	PORT MAP (Z0 => UQVN_N63, A0 => LD, A1 => UQVN_N64, A2 => D7);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N64, A0 => CS);
UQVB_B72 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N59);
UQVB_B73 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N68);
UQVB_B74 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N67);
UQVB_B75 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N66);
UQVB_B76 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N69);
UQVB_B77 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N70);
UQVB_B78 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N71);
UQVB_B79 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N65);
END lattice_arch;
-- VHDL netlist for SRRL1
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRRL1 IS 
    PORT (
        D0 : IN std_logic;
        CAIR : IN std_logic;
        CAIL : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        RL : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic
    );
END SRRL1;


ARCHITECTURE lattice_arch OF SRRL1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B2 : OR5
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => RL);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => LD);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => EN);
UQVB_B7 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N8);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => LD, A1 => UQVN_N10, A2 => D0);
UQVB_B9 : FD21
	PORT MAP (Q0 => UQVN_N8, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => EN, A1 => UQVN_N7, A2 => UQVN_N10, 
	A3 => RL, A4 => CAIR);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => EN, A1 => UQVN_N7, A2 => UQVN_N10, 
	A3 => UQVN_N1, A4 => CAIL);
END lattice_arch;
-- VHDL netlist for SRRL4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRRL4 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        CAIR : IN std_logic;
        CAIL : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        RL : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic
    );
END SRRL4;


ARCHITECTURE lattice_arch OF SRRL4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B2 : OR5
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => RL);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => LD);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => EN);
UQVB_B7 : BUF
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N8);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => LD, A1 => UQVN_N10, A2 => D0);
UQVB_B9 : FD21
	PORT MAP (Q0 => UQVN_N8, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => EN, A1 => UQVN_N7, A2 => UQVN_N10, 
	A3 => RL, A4 => CAIR);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => EN, A1 => UQVN_N7, A2 => UQVN_N10, 
	A3 => UQVN_N1, A4 => UQVN_N44);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N19, 
	A3 => UQVN_N20);
UQVB_B13 : OR5
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N12, A1 => UQVN_N13, A2 => UQVN_N14, 
	A3 => UQVN_N15, A4 => PS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => RL);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => CS);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => EN);
UQVB_B18 : BUF
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N18);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => LD, A1 => UQVN_N20, A2 => D1);
UQVB_B20 : FD21
	PORT MAP (Q0 => UQVN_N18, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B21 : AND5
	PORT MAP (Z0 => UQVN_N13, A0 => EN, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => RL, A4 => UQVN_N43);
UQVB_B22 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => EN, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => UQVN_N11, A4 => UQVN_N42);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N28, A1 => UQVN_N27, A2 => UQVN_N29, 
	A3 => UQVN_N30);
UQVB_B24 : OR5
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N22, A1 => UQVN_N23, A2 => UQVN_N24, 
	A3 => UQVN_N25, A4 => PS);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => RL);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => CS);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => LD);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => EN);
UQVB_B29 : BUF
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N28);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => LD, A1 => UQVN_N30, A2 => D2);
UQVB_B31 : FD21
	PORT MAP (Q0 => UQVN_N28, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B32 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => EN, A1 => UQVN_N27, A2 => UQVN_N30, 
	A3 => RL, A4 => UQVN_N44);
UQVB_B33 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => EN, A1 => UQVN_N27, A2 => UQVN_N30, 
	A3 => UQVN_N21, A4 => UQVN_N41);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B35 : OR5
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N33, A2 => UQVN_N34, 
	A3 => UQVN_N35, A4 => PS);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => RL);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CS);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => LD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => EN);
UQVB_B40 : BUF
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N38);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => LD, A1 => UQVN_N40, A2 => D3);
UQVB_B42 : FD21
	PORT MAP (Q0 => UQVN_N38, D0 => UQVN_N36, CLK => CLK, CD => CD);
UQVB_B43 : AND5
	PORT MAP (Z0 => UQVN_N33, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N40, 
	A3 => RL, A4 => UQVN_N42);
UQVB_B44 : AND5
	PORT MAP (Z0 => UQVN_N34, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N40, 
	A3 => UQVN_N31, A4 => CAIL);
UQVB_B45 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N43);
UQVB_B46 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N44);
UQVB_B47 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N42);
UQVB_B48 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N41);
END lattice_arch;
-- VHDL netlist for SRRL8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SRRL8 IS 
    PORT (
        D0 : IN std_logic;
        D1 : IN std_logic;
        D2 : IN std_logic;
        D3 : IN std_logic;
        D4 : IN std_logic;
        D5 : IN std_logic;
        D6 : IN std_logic;
        D7 : IN std_logic;
        CAIR : IN std_logic;
        CAIL : IN std_logic;
        CLK : IN std_logic;
        PS : IN std_logic;
        LD : IN std_logic;
        EN : IN std_logic;
        RL : IN std_logic;
        CD : IN std_logic;
        CS : IN std_logic;
        Q0 : OUT std_logic;
        Q1 : OUT std_logic;
        Q2 : OUT std_logic;
        Q3 : OUT std_logic;
        Q4 : OUT std_logic;
        Q5 : OUT std_logic;
        Q6 : OUT std_logic;
        Q7 : OUT std_logic
    );
END SRRL8;


ARCHITECTURE lattice_arch OF SRRL8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88 : std_logic;


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT BUF
    PORT (
        A0 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: BUF use  entity  lat_vhd.BUF(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT FD21
    PORT (
        D0 : IN std_logic;
        CLK : IN std_logic;
        CD : IN std_logic;
        Q0 : OUT std_logic
    );
  END COMPONENT;

for all: FD21 use  entity  lat_vhd.FD21(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


BEGIN

UQVB_B1 : AND4
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N9, 
	A3 => UQVN_N10);
UQVB_B2 : OR5
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N2, A1 => UQVN_N3, A2 => UQVN_N4, 
	A3 => UQVN_N5, A4 => PS);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => RL);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => CS);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => LD);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => EN);
UQVB_B7 : BUF
	PORT MAP (Z0 => UQVN_N84, A0 => UQVN_N8);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => LD, A1 => UQVN_N10, A2 => D0);
UQVB_B9 : FD21
	PORT MAP (Q0 => UQVN_N8, D0 => UQVN_N6, CLK => CLK, CD => CD);
UQVB_B10 : AND5
	PORT MAP (Z0 => UQVN_N3, A0 => EN, A1 => UQVN_N7, A2 => UQVN_N10, 
	A3 => RL, A4 => CAIR);
UQVB_B11 : AND5
	PORT MAP (Z0 => UQVN_N4, A0 => EN, A1 => UQVN_N7, A2 => UQVN_N10, 
	A3 => UQVN_N1, A4 => UQVN_N88);
UQVB_B12 : AND4
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N19, 
	A3 => UQVN_N20);
UQVB_B13 : OR5
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N12, A1 => UQVN_N13, A2 => UQVN_N14, 
	A3 => UQVN_N15, A4 => PS);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N11, A0 => RL);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => CS);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => LD);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => EN);
UQVB_B18 : BUF
	PORT MAP (Z0 => UQVN_N88, A0 => UQVN_N18);
UQVB_B19 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => LD, A1 => UQVN_N20, A2 => D1);
UQVB_B20 : FD21
	PORT MAP (Q0 => UQVN_N18, D0 => UQVN_N16, CLK => CLK, CD => CD);
UQVB_B21 : AND5
	PORT MAP (Z0 => UQVN_N13, A0 => EN, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => RL, A4 => UQVN_N84);
UQVB_B22 : AND5
	PORT MAP (Z0 => UQVN_N14, A0 => EN, A1 => UQVN_N17, A2 => UQVN_N20, 
	A3 => UQVN_N11, A4 => UQVN_N83);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N28, A1 => UQVN_N27, A2 => UQVN_N29, 
	A3 => UQVN_N30);
UQVB_B24 : OR5
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N22, A1 => UQVN_N23, A2 => UQVN_N24, 
	A3 => UQVN_N25, A4 => PS);
UQVB_B25 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => RL);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => CS);
UQVB_B27 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => LD);
UQVB_B28 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => EN);
UQVB_B29 : BUF
	PORT MAP (Z0 => UQVN_N83, A0 => UQVN_N28);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => LD, A1 => UQVN_N30, A2 => D2);
UQVB_B31 : FD21
	PORT MAP (Q0 => UQVN_N28, D0 => UQVN_N26, CLK => CLK, CD => CD);
UQVB_B32 : AND5
	PORT MAP (Z0 => UQVN_N23, A0 => EN, A1 => UQVN_N27, A2 => UQVN_N30, 
	A3 => RL, A4 => UQVN_N88);
UQVB_B33 : AND5
	PORT MAP (Z0 => UQVN_N24, A0 => EN, A1 => UQVN_N27, A2 => UQVN_N30, 
	A3 => UQVN_N21, A4 => UQVN_N82);
UQVB_B34 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N38, A1 => UQVN_N37, A2 => UQVN_N39, 
	A3 => UQVN_N40);
UQVB_B35 : OR5
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N32, A1 => UQVN_N33, A2 => UQVN_N34, 
	A3 => UQVN_N35, A4 => PS);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => RL);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => CS);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => LD);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => EN);
UQVB_B40 : BUF
	PORT MAP (Z0 => UQVN_N82, A0 => UQVN_N38);
UQVB_B41 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => LD, A1 => UQVN_N40, A2 => D3);
UQVB_B42 : FD21
	PORT MAP (Q0 => UQVN_N38, D0 => UQVN_N36, CLK => CLK, CD => CD);
UQVB_B43 : AND5
	PORT MAP (Z0 => UQVN_N33, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N40, 
	A3 => RL, A4 => UQVN_N83);
UQVB_B44 : AND5
	PORT MAP (Z0 => UQVN_N34, A0 => EN, A1 => UQVN_N37, A2 => UQVN_N40, 
	A3 => UQVN_N31, A4 => UQVN_N81);
UQVB_B45 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => UQVN_N48, A1 => UQVN_N47, A2 => UQVN_N49, 
	A3 => UQVN_N50);
UQVB_B46 : OR5
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N42, A1 => UQVN_N43, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => PS);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => RL);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => CS);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => LD);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => EN);
UQVB_B51 : BUF
	PORT MAP (Z0 => UQVN_N81, A0 => UQVN_N48);
UQVB_B52 : AND3
	PORT MAP (Z0 => UQVN_N45, A0 => LD, A1 => UQVN_N50, A2 => D4);
UQVB_B53 : FD21
	PORT MAP (Q0 => UQVN_N48, D0 => UQVN_N46, CLK => CLK, CD => CD);
UQVB_B54 : AND5
	PORT MAP (Z0 => UQVN_N43, A0 => EN, A1 => UQVN_N47, A2 => UQVN_N50, 
	A3 => RL, A4 => UQVN_N82);
UQVB_B55 : AND5
	PORT MAP (Z0 => UQVN_N44, A0 => EN, A1 => UQVN_N47, A2 => UQVN_N50, 
	A3 => UQVN_N41, A4 => UQVN_N87);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N58, A1 => UQVN_N57, A2 => UQVN_N59, 
	A3 => UQVN_N60);
UQVB_B57 : OR5
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N52, A1 => UQVN_N53, A2 => UQVN_N54, 
	A3 => UQVN_N55, A4 => PS);
UQVB_B58 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => RL);
UQVB_B59 : INV
	PORT MAP (ZN0 => UQVN_N60, A0 => CS);
UQVB_B60 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => LD);
UQVB_B61 : INV
	PORT MAP (ZN0 => UQVN_N59, A0 => EN);
UQVB_B62 : BUF
	PORT MAP (Z0 => UQVN_N87, A0 => UQVN_N58);
UQVB_B63 : AND3
	PORT MAP (Z0 => UQVN_N55, A0 => LD, A1 => UQVN_N60, A2 => D5);
UQVB_B64 : FD21
	PORT MAP (Q0 => UQVN_N58, D0 => UQVN_N56, CLK => CLK, CD => CD);
UQVB_B65 : AND5
	PORT MAP (Z0 => UQVN_N53, A0 => EN, A1 => UQVN_N57, A2 => UQVN_N60, 
	A3 => RL, A4 => UQVN_N81);
UQVB_B66 : AND5
	PORT MAP (Z0 => UQVN_N54, A0 => EN, A1 => UQVN_N57, A2 => UQVN_N60, 
	A3 => UQVN_N51, A4 => UQVN_N85);
UQVB_B67 : AND4
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N68, A1 => UQVN_N67, A2 => UQVN_N69, 
	A3 => UQVN_N70);
UQVB_B68 : OR5
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N62, A1 => UQVN_N63, A2 => UQVN_N64, 
	A3 => UQVN_N65, A4 => PS);
UQVB_B69 : INV
	PORT MAP (ZN0 => UQVN_N61, A0 => RL);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => CS);
UQVB_B71 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => LD);
UQVB_B72 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => EN);
UQVB_B73 : BUF
	PORT MAP (Z0 => UQVN_N85, A0 => UQVN_N68);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N65, A0 => LD, A1 => UQVN_N70, A2 => D6);
UQVB_B75 : FD21
	PORT MAP (Q0 => UQVN_N68, D0 => UQVN_N66, CLK => CLK, CD => CD);
UQVB_B76 : AND5
	PORT MAP (Z0 => UQVN_N63, A0 => EN, A1 => UQVN_N67, A2 => UQVN_N70, 
	A3 => RL, A4 => UQVN_N87);
UQVB_B77 : AND5
	PORT MAP (Z0 => UQVN_N64, A0 => EN, A1 => UQVN_N67, A2 => UQVN_N70, 
	A3 => UQVN_N61, A4 => UQVN_N86);
UQVB_B78 : AND4
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N78, A1 => UQVN_N77, A2 => UQVN_N79, 
	A3 => UQVN_N80);
UQVB_B79 : OR5
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N72, A1 => UQVN_N73, A2 => UQVN_N74, 
	A3 => UQVN_N75, A4 => PS);
UQVB_B80 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => RL);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N80, A0 => CS);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N77, A0 => LD);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N79, A0 => EN);
UQVB_B84 : BUF
	PORT MAP (Z0 => UQVN_N86, A0 => UQVN_N78);
UQVB_B85 : AND3
	PORT MAP (Z0 => UQVN_N75, A0 => LD, A1 => UQVN_N80, A2 => D7);
UQVB_B86 : FD21
	PORT MAP (Q0 => UQVN_N78, D0 => UQVN_N76, CLK => CLK, CD => CD);
UQVB_B87 : AND5
	PORT MAP (Z0 => UQVN_N73, A0 => EN, A1 => UQVN_N77, A2 => UQVN_N80, 
	A3 => RL, A4 => UQVN_N85);
UQVB_B88 : AND5
	PORT MAP (Z0 => UQVN_N74, A0 => EN, A1 => UQVN_N77, A2 => UQVN_N80, 
	A3 => UQVN_N71, A4 => CAIL);
UQVB_B89 : BUF
	PORT MAP (Z0 => Q7, A0 => UQVN_N86);
UQVB_B90 : BUF
	PORT MAP (Z0 => Q6, A0 => UQVN_N85);
UQVB_B91 : BUF
	PORT MAP (Z0 => Q4, A0 => UQVN_N81);
UQVB_B92 : BUF
	PORT MAP (Z0 => Q5, A0 => UQVN_N87);
UQVB_B93 : BUF
	PORT MAP (Z0 => Q0, A0 => UQVN_N84);
UQVB_B94 : BUF
	PORT MAP (Z0 => Q1, A0 => UQVN_N88);
UQVB_B95 : BUF
	PORT MAP (Z0 => Q3, A0 => UQVN_N82);
UQVB_B96 : BUF
	PORT MAP (Z0 => Q2, A0 => UQVN_N83);
END lattice_arch;
-- VHDL netlist for SUBF1
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBF1 IS 
    PORT (
        A0 : IN std_logic;
        B0 : IN std_logic;
        BI : IN std_logic;
        Z0 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBF1;


ARCHITECTURE lattice_arch OF SUBF1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9 : std_logic;


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


BEGIN

UQVB_B1 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N4);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N9, A1 => BI);
UQVB_B3 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => B0, A1 => UQVN_N1);
UQVB_B4 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => A0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => B0);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => BI);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => BI, A1 => B0);
UQVB_B9 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => BI, A1 => UQVN_N5);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N8, A0 => B0, A1 => UQVN_N5);
UQVB_B11 : OR3
	PORT MAP (Z0 => BO, A0 => UQVN_N6, A1 => UQVN_N7, A2 => UQVN_N8);
END lattice_arch;
-- VHDL netlist for SUBF16A
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBF16A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B10 : IN std_logic;
        B11 : IN std_logic;
        B12 : IN std_logic;
        B13 : IN std_logic;
        B14 : IN std_logic;
        B15 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        B8 : IN std_logic;
        B9 : IN std_logic;
        BI : IN std_logic;
        BO : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z10 : OUT std_logic;
        Z11 : OUT std_logic;
        Z12 : OUT std_logic;
        Z13 : OUT std_logic;
        Z14 : OUT std_logic;
        Z15 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        Z8 : OUT std_logic;
        Z9 : OUT std_logic
    );
END SUBF16A;


ARCHITECTURE lattice_arch OF SUBF16A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 UQVN_N113, UQVN_N114, UQVN_N115, UQVN_N116,
	 UQVN_N117, UQVN_N118, UQVN_N119, UQVN_N120,
	 UQVN_N121, UQVN_N122, UQVN_N123, UQVN_N124,
	 UQVN_N125, UQVN_N126, UQVN_N127, UQVN_N128,
	 UQVN_N129, UQVN_N130, UQVN_N131, UQVN_N132,
	 UQVN_N133, UQVN_N134, UQVN_N135, UQVN_N136,
	 UQVN_N137, UQVN_N138, UQVN_N139, UQVN_N140,
	 UQVN_N141, UQVN_N142, UQVN_N143, UQVN_N144,
	 UQVN_N145, UQVN_N146, UQVN_N147, UQVN_N148,
	 UQVN_N149, UQVN_N150, UQVN_N151, UQVN_N152,
	 UQVN_N153, UQVN_N154, UQVN_N155, UQVN_N156,
	 UQVN_N157, UQVN_N158, UQVN_N159, UQVN_N160,
	 UQVN_N161, UQVN_N162, UQVN_N163, UQVN_N164,
	 UQVN_N165, UQVN_N166, UQVN_N167, UQVN_N168,
	 UQVN_N169, UQVN_N170, UQVN_N171, UQVN_N172,
	 UQVN_N173, UQVN_N174, UQVN_N175, UQVN_N176,
	 UQVN_N177, UQVN_N178, UQVN_N179, UQVN_N180,
	 UQVN_N181, UQVN_N182, UQVN_N183, UQVN_N184,
	 UQVN_N185, UQVN_N186, UQVN_N187, UQVN_N188,
	 UQVN_N189, UQVN_N190, UQVN_N191, UQVN_N192,
	 UQVN_N193, UQVN_N194, UQVN_N195, UQVN_N196,
	 UQVN_N197, UQVN_N198, UQVN_N199, UQVN_N200,
	 UQVN_N201, UQVN_N202, UQVN_N203, UQVN_N204,
	 UQVN_N205, UQVN_N206, UQVN_N207, UQVN_N208,
	 UQVN_N209, UQVN_N210, UQVN_N211, UQVN_N212,
	 UQVN_N213, UQVN_N214, UQVN_N215, UQVN_N216,
	 UQVN_N217, UQVN_N218, UQVN_N219, UQVN_N220,
	 UQVN_N221, UQVN_N222, UQVN_N223, UQVN_N224,
	 UQVN_N225, UQVN_N226, UQVN_N227, UQVN_N228,
	 UQVN_N229, UQVN_N230, UQVN_N231, UQVN_N232,
	 UQVN_N233, UQVN_N234, UQVN_N235, UQVN_N236,
	 UQVN_N237, UQVN_N238, UQVN_N239, UQVN_N240,
	 G012, G1214, G345, G678,
	 G911, P012, P1214, P345,
	 P678, P911 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => P345, A1 => UQVN_N240);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N236, A0 => G345, A1 => UQVN_N1);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N237, A0 => G678, A1 => UQVN_N2, A2 => UQVN_N3);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => P678, A1 => P345, A2 => UQVN_N240);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => P678, A1 => G345);
UQVB_B6 : OR4
	PORT MAP (Z0 => UQVN_N238, A0 => G911, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => UQVN_N6);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => P911, A1 => G678);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => P911, A1 => P678, A2 => G345);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => P911, A1 => P678, A2 => P345, 
	A3 => UQVN_N240);
UQVB_B10 : OR5
	PORT MAP (Z0 => UQVN_N239, A0 => G1214, A1 => UQVN_N7, A2 => UQVN_N8, 
	A3 => UQVN_N9, A4 => UQVN_N10);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => P1214, A1 => G911);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => P1214, A1 => P911, A2 => G678);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => G345);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => P345, A4 => UQVN_N240);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => P012, A1 => BI);
UQVB_B16 : OR2
	PORT MAP (Z0 => UQVN_N240, A0 => G012, A1 => UQVN_N11);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => BI);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => B1);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => B2);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => A0);
UQVB_B21 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N51, A1 => BI);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N13, A0 => B0, A1 => UQVN_N54);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N12, A1 => UQVN_N13);
UQVB_B24 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N14);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => A0, A1 => B1, A2 => UQVN_N51);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N52, A1 => B0, A2 => BI);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N48, A1 => UQVN_N52, A2 => BI);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => B1, A1 => UQVN_N51, A2 => UQVN_N54);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => A0, A1 => B1, A2 => UQVN_N54);
UQVB_B30 : OR6
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N15, 
	A3 => UQVN_N16, A4 => UQVN_N20, A5 => UQVN_N19);
UQVB_B31 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N21);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N48, A1 => UQVN_N52, A2 => B0);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N48, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B34 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N49, A1 => B1, A2 => B2);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N48, A1 => UQVN_N50, A2 => B0, 
	A3 => B1);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N50, A1 => B2);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N48, A1 => UQVN_N49, A2 => B0, 
	A3 => B2);
UQVB_B38 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N49, A1 => UQVN_N50, A2 => B1);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N48, A1 => UQVN_N49, A2 => UQVN_N50, 
	A3 => B0);
UQVB_B40 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N22, A4 => UQVN_N26, A5 => UQVN_N27, A6 => UQVN_N28);
UQVB_B41 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => A0, A1 => UQVN_N51);
UQVB_B42 : AND2
	PORT MAP (Z0 => UQVN_N29, A0 => A1, A1 => UQVN_N52);
UQVB_B43 : AND2
	PORT MAP (Z0 => UQVN_N30, A0 => A2, A1 => UQVN_N53);
UQVB_B44 : NOR3
	PORT MAP (ZN0 => P012, A0 => UQVN_N31, A1 => UQVN_N29, A2 => UQVN_N30);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => B0);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => A1);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => A2);
UQVB_B48 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N45);
UQVB_B49 : AND4
	PORT MAP (Z0 => UQVN_N44, A0 => A0, A1 => A1, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B50 : AND4
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N48, A1 => UQVN_N49, A2 => UQVN_N53, 
	A3 => BI);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N43, A0 => A0, A1 => A1, A2 => UQVN_N51, 
	A3 => B2);
UQVB_B52 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => A1, A1 => UQVN_N51, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B53 : AND4
	PORT MAP (Z0 => UQVN_N41, A0 => UQVN_N48, A1 => UQVN_N49, A2 => B0, 
	A3 => UQVN_N53);
UQVB_B54 : AND4
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N49, A1 => B0, A2 => UQVN_N53, 
	A3 => BI);
UQVB_B55 : AND4
	PORT MAP (Z0 => UQVN_N39, A0 => A0, A1 => UQVN_N52, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B56 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => A0, A1 => UQVN_N51, A2 => UQVN_N52, 
	A3 => B2);
UQVB_B57 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N51, A1 => UQVN_N52, A2 => B2, 
	A3 => UQVN_N54);
UQVB_B58 : AND3
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N49, A1 => UQVN_N53, A2 => B1);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N48, A1 => B1, A2 => UQVN_N53, 
	A3 => BI);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N48, A1 => B0, A2 => B1, 
	A3 => UQVN_N53);
UQVB_B61 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => A1, A1 => UQVN_N52, A2 => B2);
UQVB_B62 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => B0, A1 => B1, A2 => UQVN_N53, 
	A3 => BI);
UQVB_B63 : OR12
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N43, A1 => UQVN_N42, A2 => UQVN_N41, 
	A3 => UQVN_N40, A4 => UQVN_N39, A5 => UQVN_N38, A6 => UQVN_N37, 
	A7 => UQVN_N36, A8 => UQVN_N35, A9 => UQVN_N34, A10 => UQVN_N33, 
	A11 => UQVN_N32);
UQVB_B64 : OR3
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N44, A1 => UQVN_N46, A2 => UQVN_N47);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N97, A0 => UQVN_N240);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N95, A0 => B4);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N96, A0 => B5);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N91, A0 => A3);
UQVB_B69 : AND2
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N94, A1 => UQVN_N240);
UQVB_B70 : AND2
	PORT MAP (Z0 => UQVN_N56, A0 => B3, A1 => UQVN_N97);
UQVB_B71 : OR2
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N55, A1 => UQVN_N56);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N57);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N63, A0 => A3, A1 => B4, A2 => UQVN_N94);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N95, A1 => B3, A2 => UQVN_N240);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N91, A1 => UQVN_N95, A2 => UQVN_N240);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N60, A0 => B4, A1 => UQVN_N94, A2 => UQVN_N97);
UQVB_B77 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => A3, A1 => B4, A2 => UQVN_N97);
UQVB_B78 : OR6
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N61, A1 => UQVN_N60, A2 => UQVN_N58, 
	A3 => UQVN_N59, A4 => UQVN_N63, A5 => UQVN_N62);
UQVB_B79 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N64);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N91, A1 => UQVN_N95, A2 => B3);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N68, A0 => UQVN_N91, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B82 : AND3
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N92, A1 => B4, A2 => B5);
UQVB_B83 : AND4
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N91, A1 => UQVN_N93, A2 => B3, 
	A3 => B4);
UQVB_B84 : AND2
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N93, A1 => B5);
UQVB_B85 : AND4
	PORT MAP (Z0 => UQVN_N69, A0 => UQVN_N91, A1 => UQVN_N92, A2 => B3, 
	A3 => B5);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N92, A1 => UQVN_N93, A2 => B4);
UQVB_B87 : AND4
	PORT MAP (Z0 => UQVN_N71, A0 => UQVN_N91, A1 => UQVN_N92, A2 => UQVN_N93, 
	A3 => B3);
UQVB_B88 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N68, A1 => UQVN_N67, A2 => UQVN_N66, 
	A3 => UQVN_N65, A4 => UQVN_N69, A5 => UQVN_N70, A6 => UQVN_N71);
UQVB_B89 : AND2
	PORT MAP (Z0 => UQVN_N74, A0 => A3, A1 => UQVN_N94);
UQVB_B90 : AND2
	PORT MAP (Z0 => UQVN_N72, A0 => A4, A1 => UQVN_N95);
UQVB_B91 : AND2
	PORT MAP (Z0 => UQVN_N73, A0 => A5, A1 => UQVN_N96);
UQVB_B92 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N74, A1 => UQVN_N72, A2 => UQVN_N73);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N94, A0 => B3);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N92, A0 => A4);
UQVB_B95 : INV
	PORT MAP (ZN0 => UQVN_N93, A0 => A5);
UQVB_B96 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N88);
UQVB_B97 : AND4
	PORT MAP (Z0 => UQVN_N87, A0 => A3, A1 => A4, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B98 : AND4
	PORT MAP (Z0 => UQVN_N89, A0 => UQVN_N91, A1 => UQVN_N92, A2 => UQVN_N96, 
	A3 => UQVN_N240);
UQVB_B99 : AND4
	PORT MAP (Z0 => UQVN_N86, A0 => A3, A1 => A4, A2 => UQVN_N94, 
	A3 => B5);
UQVB_B100 : AND4
	PORT MAP (Z0 => UQVN_N85, A0 => A4, A1 => UQVN_N94, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B101 : AND4
	PORT MAP (Z0 => UQVN_N84, A0 => UQVN_N91, A1 => UQVN_N92, A2 => B3, 
	A3 => UQVN_N96);
UQVB_B102 : AND4
	PORT MAP (Z0 => UQVN_N83, A0 => UQVN_N92, A1 => B3, A2 => UQVN_N96, 
	A3 => UQVN_N240);
UQVB_B103 : AND4
	PORT MAP (Z0 => UQVN_N82, A0 => A3, A1 => UQVN_N95, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B104 : AND4
	PORT MAP (Z0 => UQVN_N81, A0 => A3, A1 => UQVN_N94, A2 => UQVN_N95, 
	A3 => B5);
UQVB_B105 : AND4
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N94, A1 => UQVN_N95, A2 => B5, 
	A3 => UQVN_N97);
UQVB_B106 : AND3
	PORT MAP (Z0 => UQVN_N79, A0 => UQVN_N92, A1 => UQVN_N96, A2 => B4);
UQVB_B107 : AND4
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N91, A1 => B4, A2 => UQVN_N96, 
	A3 => UQVN_N240);
UQVB_B108 : AND4
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N91, A1 => B3, A2 => B4, 
	A3 => UQVN_N96);
UQVB_B109 : AND3
	PORT MAP (Z0 => UQVN_N76, A0 => A4, A1 => UQVN_N95, A2 => B5);
UQVB_B110 : AND4
	PORT MAP (Z0 => UQVN_N75, A0 => B3, A1 => B4, A2 => UQVN_N96, 
	A3 => UQVN_N240);
UQVB_B111 : OR12
	PORT MAP (Z0 => UQVN_N90, A0 => UQVN_N86, A1 => UQVN_N85, A2 => UQVN_N84, 
	A3 => UQVN_N83, A4 => UQVN_N82, A5 => UQVN_N81, A6 => UQVN_N80, 
	A7 => UQVN_N79, A8 => UQVN_N78, A9 => UQVN_N77, A10 => UQVN_N76, 
	A11 => UQVN_N75);
UQVB_B112 : OR3
	PORT MAP (Z0 => UQVN_N88, A0 => UQVN_N87, A1 => UQVN_N89, A2 => UQVN_N90);
UQVB_B113 : INV
	PORT MAP (ZN0 => UQVN_N140, A0 => UQVN_N236);
UQVB_B114 : INV
	PORT MAP (ZN0 => UQVN_N138, A0 => B7);
UQVB_B115 : INV
	PORT MAP (ZN0 => UQVN_N139, A0 => B8);
UQVB_B116 : INV
	PORT MAP (ZN0 => UQVN_N134, A0 => A6);
UQVB_B117 : AND2
	PORT MAP (Z0 => UQVN_N98, A0 => UQVN_N137, A1 => UQVN_N236);
UQVB_B118 : AND2
	PORT MAP (Z0 => UQVN_N99, A0 => B6, A1 => UQVN_N140);
UQVB_B119 : OR2
	PORT MAP (Z0 => UQVN_N100, A0 => UQVN_N98, A1 => UQVN_N99);
UQVB_B120 : LXOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N100);
UQVB_B121 : AND3
	PORT MAP (Z0 => UQVN_N106, A0 => A6, A1 => B7, A2 => UQVN_N137);
UQVB_B122 : AND3
	PORT MAP (Z0 => UQVN_N102, A0 => UQVN_N138, A1 => B6, A2 => UQVN_N236);
UQVB_B123 : AND3
	PORT MAP (Z0 => UQVN_N101, A0 => UQVN_N134, A1 => UQVN_N138, A2 => UQVN_N236);
UQVB_B124 : AND3
	PORT MAP (Z0 => UQVN_N103, A0 => B7, A1 => UQVN_N137, A2 => UQVN_N140);
UQVB_B125 : AND3
	PORT MAP (Z0 => UQVN_N104, A0 => A6, A1 => B7, A2 => UQVN_N140);
UQVB_B126 : OR6
	PORT MAP (Z0 => UQVN_N107, A0 => UQVN_N104, A1 => UQVN_N103, A2 => UQVN_N101, 
	A3 => UQVN_N102, A4 => UQVN_N106, A5 => UQVN_N105);
UQVB_B127 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N107);
UQVB_B128 : AND3
	PORT MAP (Z0 => UQVN_N105, A0 => UQVN_N134, A1 => UQVN_N138, A2 => B6);
UQVB_B129 : AND4
	PORT MAP (Z0 => UQVN_N111, A0 => UQVN_N134, A1 => B6, A2 => B7, 
	A3 => B8);
UQVB_B130 : AND3
	PORT MAP (Z0 => UQVN_N110, A0 => UQVN_N135, A1 => B7, A2 => B8);
UQVB_B131 : AND4
	PORT MAP (Z0 => UQVN_N109, A0 => UQVN_N134, A1 => UQVN_N136, A2 => B6, 
	A3 => B7);
UQVB_B132 : AND2
	PORT MAP (Z0 => UQVN_N108, A0 => UQVN_N136, A1 => B8);
UQVB_B133 : AND4
	PORT MAP (Z0 => UQVN_N112, A0 => UQVN_N134, A1 => UQVN_N135, A2 => B6, 
	A3 => B8);
UQVB_B134 : AND3
	PORT MAP (Z0 => UQVN_N113, A0 => UQVN_N135, A1 => UQVN_N136, A2 => B7);
UQVB_B135 : AND4
	PORT MAP (Z0 => UQVN_N114, A0 => UQVN_N134, A1 => UQVN_N135, A2 => UQVN_N136, 
	A3 => B6);
UQVB_B136 : OR7
	PORT MAP (Z0 => G678, A0 => UQVN_N111, A1 => UQVN_N110, A2 => UQVN_N109, 
	A3 => UQVN_N108, A4 => UQVN_N112, A5 => UQVN_N113, A6 => UQVN_N114);
UQVB_B137 : AND2
	PORT MAP (Z0 => UQVN_N117, A0 => A6, A1 => UQVN_N137);
UQVB_B138 : AND2
	PORT MAP (Z0 => UQVN_N115, A0 => A7, A1 => UQVN_N138);
UQVB_B139 : AND2
	PORT MAP (Z0 => UQVN_N116, A0 => A8, A1 => UQVN_N139);
UQVB_B140 : NOR3
	PORT MAP (ZN0 => P678, A0 => UQVN_N117, A1 => UQVN_N115, A2 => UQVN_N116);
UQVB_B141 : INV
	PORT MAP (ZN0 => UQVN_N137, A0 => B6);
UQVB_B142 : INV
	PORT MAP (ZN0 => UQVN_N135, A0 => A7);
UQVB_B143 : INV
	PORT MAP (ZN0 => UQVN_N136, A0 => A8);
UQVB_B144 : LXOR2
	PORT MAP (Z0 => Z8, A0 => A8, A1 => UQVN_N131);
UQVB_B145 : AND4
	PORT MAP (Z0 => UQVN_N130, A0 => A6, A1 => A7, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B146 : AND4
	PORT MAP (Z0 => UQVN_N132, A0 => UQVN_N134, A1 => UQVN_N135, A2 => UQVN_N139, 
	A3 => UQVN_N236);
UQVB_B147 : AND4
	PORT MAP (Z0 => UQVN_N129, A0 => A6, A1 => A7, A2 => UQVN_N137, 
	A3 => B8);
UQVB_B148 : AND4
	PORT MAP (Z0 => UQVN_N128, A0 => A7, A1 => UQVN_N137, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B149 : AND4
	PORT MAP (Z0 => UQVN_N127, A0 => UQVN_N134, A1 => UQVN_N135, A2 => B6, 
	A3 => UQVN_N139);
UQVB_B150 : AND4
	PORT MAP (Z0 => UQVN_N126, A0 => UQVN_N135, A1 => B6, A2 => UQVN_N139, 
	A3 => UQVN_N236);
UQVB_B151 : AND4
	PORT MAP (Z0 => UQVN_N125, A0 => A6, A1 => UQVN_N138, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B152 : AND4
	PORT MAP (Z0 => UQVN_N124, A0 => A6, A1 => UQVN_N137, A2 => UQVN_N138, 
	A3 => B8);
UQVB_B153 : AND4
	PORT MAP (Z0 => UQVN_N123, A0 => UQVN_N137, A1 => UQVN_N138, A2 => B8, 
	A3 => UQVN_N140);
UQVB_B154 : AND3
	PORT MAP (Z0 => UQVN_N122, A0 => UQVN_N135, A1 => UQVN_N139, A2 => B7);
UQVB_B155 : AND4
	PORT MAP (Z0 => UQVN_N121, A0 => UQVN_N134, A1 => B7, A2 => UQVN_N139, 
	A3 => UQVN_N236);
UQVB_B156 : AND4
	PORT MAP (Z0 => UQVN_N120, A0 => UQVN_N134, A1 => B6, A2 => B7, 
	A3 => UQVN_N139);
UQVB_B157 : AND3
	PORT MAP (Z0 => UQVN_N119, A0 => A7, A1 => UQVN_N138, A2 => B8);
UQVB_B158 : AND4
	PORT MAP (Z0 => UQVN_N118, A0 => B6, A1 => B7, A2 => UQVN_N139, 
	A3 => UQVN_N236);
UQVB_B159 : OR12
	PORT MAP (Z0 => UQVN_N133, A0 => UQVN_N129, A1 => UQVN_N128, A2 => UQVN_N127, 
	A3 => UQVN_N126, A4 => UQVN_N125, A5 => UQVN_N124, A6 => UQVN_N123, 
	A7 => UQVN_N122, A8 => UQVN_N121, A9 => UQVN_N120, A10 => UQVN_N119, 
	A11 => UQVN_N118);
UQVB_B160 : OR3
	PORT MAP (Z0 => UQVN_N131, A0 => UQVN_N130, A1 => UQVN_N132, A2 => UQVN_N133);
UQVB_B161 : INV
	PORT MAP (ZN0 => UQVN_N183, A0 => UQVN_N237);
UQVB_B162 : INV
	PORT MAP (ZN0 => UQVN_N181, A0 => B10);
UQVB_B163 : INV
	PORT MAP (ZN0 => UQVN_N182, A0 => B11);
UQVB_B164 : INV
	PORT MAP (ZN0 => UQVN_N177, A0 => A9);
UQVB_B165 : AND2
	PORT MAP (Z0 => UQVN_N141, A0 => UQVN_N180, A1 => UQVN_N237);
UQVB_B166 : AND2
	PORT MAP (Z0 => UQVN_N142, A0 => B9, A1 => UQVN_N183);
UQVB_B167 : OR2
	PORT MAP (Z0 => UQVN_N143, A0 => UQVN_N141, A1 => UQVN_N142);
UQVB_B168 : LXOR2
	PORT MAP (Z0 => Z9, A0 => A9, A1 => UQVN_N143);
UQVB_B169 : AND3
	PORT MAP (Z0 => UQVN_N149, A0 => A9, A1 => B10, A2 => UQVN_N180);
UQVB_B170 : AND3
	PORT MAP (Z0 => UQVN_N145, A0 => UQVN_N181, A1 => B9, A2 => UQVN_N237);
UQVB_B171 : AND3
	PORT MAP (Z0 => UQVN_N144, A0 => UQVN_N177, A1 => UQVN_N181, A2 => UQVN_N237);
UQVB_B172 : AND3
	PORT MAP (Z0 => UQVN_N146, A0 => B10, A1 => UQVN_N180, A2 => UQVN_N183);
UQVB_B173 : AND3
	PORT MAP (Z0 => UQVN_N147, A0 => A9, A1 => B10, A2 => UQVN_N183);
UQVB_B174 : OR6
	PORT MAP (Z0 => UQVN_N150, A0 => UQVN_N147, A1 => UQVN_N146, A2 => UQVN_N144, 
	A3 => UQVN_N145, A4 => UQVN_N149, A5 => UQVN_N148);
UQVB_B175 : LXOR2
	PORT MAP (Z0 => Z10, A0 => A10, A1 => UQVN_N150);
UQVB_B176 : AND3
	PORT MAP (Z0 => UQVN_N148, A0 => UQVN_N177, A1 => UQVN_N181, A2 => B9);
UQVB_B177 : AND4
	PORT MAP (Z0 => UQVN_N154, A0 => UQVN_N177, A1 => B9, A2 => B10, 
	A3 => B11);
UQVB_B178 : AND3
	PORT MAP (Z0 => UQVN_N153, A0 => UQVN_N178, A1 => B10, A2 => B11);
UQVB_B179 : AND4
	PORT MAP (Z0 => UQVN_N152, A0 => UQVN_N177, A1 => UQVN_N179, A2 => B9, 
	A3 => B10);
UQVB_B180 : AND2
	PORT MAP (Z0 => UQVN_N151, A0 => UQVN_N179, A1 => B11);
UQVB_B181 : AND4
	PORT MAP (Z0 => UQVN_N155, A0 => UQVN_N177, A1 => UQVN_N178, A2 => B9, 
	A3 => B11);
UQVB_B182 : AND3
	PORT MAP (Z0 => UQVN_N156, A0 => UQVN_N178, A1 => UQVN_N179, A2 => B10);
UQVB_B183 : AND4
	PORT MAP (Z0 => UQVN_N157, A0 => UQVN_N177, A1 => UQVN_N178, A2 => UQVN_N179, 
	A3 => B9);
UQVB_B184 : OR7
	PORT MAP (Z0 => G911, A0 => UQVN_N154, A1 => UQVN_N153, A2 => UQVN_N152, 
	A3 => UQVN_N151, A4 => UQVN_N155, A5 => UQVN_N156, A6 => UQVN_N157);
UQVB_B185 : AND2
	PORT MAP (Z0 => UQVN_N160, A0 => A9, A1 => UQVN_N180);
UQVB_B186 : AND2
	PORT MAP (Z0 => UQVN_N158, A0 => A10, A1 => UQVN_N181);
UQVB_B187 : AND2
	PORT MAP (Z0 => UQVN_N159, A0 => A11, A1 => UQVN_N182);
UQVB_B188 : NOR3
	PORT MAP (ZN0 => P911, A0 => UQVN_N160, A1 => UQVN_N158, A2 => UQVN_N159);
UQVB_B189 : INV
	PORT MAP (ZN0 => UQVN_N180, A0 => B9);
UQVB_B190 : INV
	PORT MAP (ZN0 => UQVN_N178, A0 => A10);
UQVB_B191 : INV
	PORT MAP (ZN0 => UQVN_N179, A0 => A11);
UQVB_B192 : LXOR2
	PORT MAP (Z0 => Z11, A0 => A11, A1 => UQVN_N174);
UQVB_B193 : AND4
	PORT MAP (Z0 => UQVN_N173, A0 => A9, A1 => A10, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B194 : AND4
	PORT MAP (Z0 => UQVN_N175, A0 => UQVN_N177, A1 => UQVN_N178, A2 => UQVN_N182, 
	A3 => UQVN_N237);
UQVB_B195 : AND4
	PORT MAP (Z0 => UQVN_N172, A0 => A9, A1 => A10, A2 => UQVN_N180, 
	A3 => B11);
UQVB_B196 : AND4
	PORT MAP (Z0 => UQVN_N171, A0 => A10, A1 => UQVN_N180, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B197 : AND4
	PORT MAP (Z0 => UQVN_N170, A0 => UQVN_N177, A1 => UQVN_N178, A2 => B9, 
	A3 => UQVN_N182);
UQVB_B198 : AND4
	PORT MAP (Z0 => UQVN_N169, A0 => UQVN_N178, A1 => B9, A2 => UQVN_N182, 
	A3 => UQVN_N237);
UQVB_B199 : AND4
	PORT MAP (Z0 => UQVN_N168, A0 => A9, A1 => UQVN_N181, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B200 : AND4
	PORT MAP (Z0 => UQVN_N167, A0 => A9, A1 => UQVN_N180, A2 => UQVN_N181, 
	A3 => B11);
UQVB_B201 : AND4
	PORT MAP (Z0 => UQVN_N166, A0 => UQVN_N180, A1 => UQVN_N181, A2 => B11, 
	A3 => UQVN_N183);
UQVB_B202 : AND3
	PORT MAP (Z0 => UQVN_N165, A0 => UQVN_N178, A1 => UQVN_N182, A2 => B10);
UQVB_B203 : AND4
	PORT MAP (Z0 => UQVN_N164, A0 => UQVN_N177, A1 => B10, A2 => UQVN_N182, 
	A3 => UQVN_N237);
UQVB_B204 : AND4
	PORT MAP (Z0 => UQVN_N163, A0 => UQVN_N177, A1 => B9, A2 => B10, 
	A3 => UQVN_N182);
UQVB_B205 : AND3
	PORT MAP (Z0 => UQVN_N162, A0 => A10, A1 => UQVN_N181, A2 => B11);
UQVB_B206 : AND4
	PORT MAP (Z0 => UQVN_N161, A0 => B9, A1 => B10, A2 => UQVN_N182, 
	A3 => UQVN_N237);
UQVB_B207 : OR12
	PORT MAP (Z0 => UQVN_N176, A0 => UQVN_N172, A1 => UQVN_N171, A2 => UQVN_N170, 
	A3 => UQVN_N169, A4 => UQVN_N168, A5 => UQVN_N167, A6 => UQVN_N166, 
	A7 => UQVN_N165, A8 => UQVN_N164, A9 => UQVN_N163, A10 => UQVN_N162, 
	A11 => UQVN_N161);
UQVB_B208 : OR3
	PORT MAP (Z0 => UQVN_N174, A0 => UQVN_N173, A1 => UQVN_N175, A2 => UQVN_N176);
UQVB_B209 : INV
	PORT MAP (ZN0 => UQVN_N226, A0 => UQVN_N238);
UQVB_B210 : INV
	PORT MAP (ZN0 => UQVN_N224, A0 => B13);
UQVB_B211 : INV
	PORT MAP (ZN0 => UQVN_N225, A0 => B14);
UQVB_B212 : INV
	PORT MAP (ZN0 => UQVN_N220, A0 => A12);
UQVB_B213 : AND2
	PORT MAP (Z0 => UQVN_N184, A0 => UQVN_N223, A1 => UQVN_N238);
UQVB_B214 : AND2
	PORT MAP (Z0 => UQVN_N185, A0 => B12, A1 => UQVN_N226);
UQVB_B215 : OR2
	PORT MAP (Z0 => UQVN_N186, A0 => UQVN_N184, A1 => UQVN_N185);
UQVB_B216 : LXOR2
	PORT MAP (Z0 => Z12, A0 => A12, A1 => UQVN_N186);
UQVB_B217 : AND3
	PORT MAP (Z0 => UQVN_N192, A0 => A12, A1 => B13, A2 => UQVN_N223);
UQVB_B218 : AND3
	PORT MAP (Z0 => UQVN_N188, A0 => UQVN_N224, A1 => B12, A2 => UQVN_N238);
UQVB_B219 : AND3
	PORT MAP (Z0 => UQVN_N187, A0 => UQVN_N220, A1 => UQVN_N224, A2 => UQVN_N238);
UQVB_B220 : AND3
	PORT MAP (Z0 => UQVN_N189, A0 => B13, A1 => UQVN_N223, A2 => UQVN_N226);
UQVB_B221 : AND3
	PORT MAP (Z0 => UQVN_N190, A0 => A12, A1 => B13, A2 => UQVN_N226);
UQVB_B222 : OR6
	PORT MAP (Z0 => UQVN_N193, A0 => UQVN_N190, A1 => UQVN_N189, A2 => UQVN_N187, 
	A3 => UQVN_N188, A4 => UQVN_N192, A5 => UQVN_N191);
UQVB_B223 : LXOR2
	PORT MAP (Z0 => Z13, A0 => A13, A1 => UQVN_N193);
UQVB_B224 : AND3
	PORT MAP (Z0 => UQVN_N191, A0 => UQVN_N220, A1 => UQVN_N224, A2 => B12);
UQVB_B225 : AND4
	PORT MAP (Z0 => UQVN_N197, A0 => UQVN_N220, A1 => B12, A2 => B13, 
	A3 => B14);
UQVB_B226 : AND3
	PORT MAP (Z0 => UQVN_N196, A0 => UQVN_N221, A1 => B13, A2 => B14);
UQVB_B227 : AND4
	PORT MAP (Z0 => UQVN_N195, A0 => UQVN_N220, A1 => UQVN_N222, A2 => B12, 
	A3 => B13);
UQVB_B228 : AND2
	PORT MAP (Z0 => UQVN_N194, A0 => UQVN_N222, A1 => B14);
UQVB_B229 : AND4
	PORT MAP (Z0 => UQVN_N198, A0 => UQVN_N220, A1 => UQVN_N221, A2 => B12, 
	A3 => B14);
UQVB_B230 : AND3
	PORT MAP (Z0 => UQVN_N199, A0 => UQVN_N221, A1 => UQVN_N222, A2 => B13);
UQVB_B231 : AND4
	PORT MAP (Z0 => UQVN_N200, A0 => UQVN_N220, A1 => UQVN_N221, A2 => UQVN_N222, 
	A3 => B12);
UQVB_B232 : OR7
	PORT MAP (Z0 => G1214, A0 => UQVN_N197, A1 => UQVN_N196, A2 => UQVN_N195, 
	A3 => UQVN_N194, A4 => UQVN_N198, A5 => UQVN_N199, A6 => UQVN_N200);
UQVB_B233 : AND2
	PORT MAP (Z0 => UQVN_N203, A0 => A12, A1 => UQVN_N223);
UQVB_B234 : AND2
	PORT MAP (Z0 => UQVN_N201, A0 => A13, A1 => UQVN_N224);
UQVB_B235 : AND2
	PORT MAP (Z0 => UQVN_N202, A0 => A14, A1 => UQVN_N225);
UQVB_B236 : NOR3
	PORT MAP (ZN0 => P1214, A0 => UQVN_N203, A1 => UQVN_N201, A2 => UQVN_N202);
UQVB_B237 : INV
	PORT MAP (ZN0 => UQVN_N223, A0 => B12);
UQVB_B238 : INV
	PORT MAP (ZN0 => UQVN_N221, A0 => A13);
UQVB_B239 : INV
	PORT MAP (ZN0 => UQVN_N222, A0 => A14);
UQVB_B240 : LXOR2
	PORT MAP (Z0 => Z14, A0 => A14, A1 => UQVN_N217);
UQVB_B241 : AND4
	PORT MAP (Z0 => UQVN_N216, A0 => A12, A1 => A13, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B242 : AND4
	PORT MAP (Z0 => UQVN_N218, A0 => UQVN_N220, A1 => UQVN_N221, A2 => UQVN_N225, 
	A3 => UQVN_N238);
UQVB_B243 : AND4
	PORT MAP (Z0 => UQVN_N215, A0 => A12, A1 => A13, A2 => UQVN_N223, 
	A3 => B14);
UQVB_B244 : AND4
	PORT MAP (Z0 => UQVN_N214, A0 => A13, A1 => UQVN_N223, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B245 : AND4
	PORT MAP (Z0 => UQVN_N213, A0 => UQVN_N220, A1 => UQVN_N221, A2 => B12, 
	A3 => UQVN_N225);
UQVB_B246 : AND4
	PORT MAP (Z0 => UQVN_N212, A0 => UQVN_N221, A1 => B12, A2 => UQVN_N225, 
	A3 => UQVN_N238);
UQVB_B247 : AND4
	PORT MAP (Z0 => UQVN_N211, A0 => A12, A1 => UQVN_N224, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B248 : AND4
	PORT MAP (Z0 => UQVN_N210, A0 => A12, A1 => UQVN_N223, A2 => UQVN_N224, 
	A3 => B14);
UQVB_B249 : AND4
	PORT MAP (Z0 => UQVN_N209, A0 => UQVN_N223, A1 => UQVN_N224, A2 => B14, 
	A3 => UQVN_N226);
UQVB_B250 : AND3
	PORT MAP (Z0 => UQVN_N208, A0 => UQVN_N221, A1 => UQVN_N225, A2 => B13);
UQVB_B251 : AND4
	PORT MAP (Z0 => UQVN_N207, A0 => UQVN_N220, A1 => B13, A2 => UQVN_N225, 
	A3 => UQVN_N238);
UQVB_B252 : AND4
	PORT MAP (Z0 => UQVN_N206, A0 => UQVN_N220, A1 => B12, A2 => B13, 
	A3 => UQVN_N225);
UQVB_B253 : AND3
	PORT MAP (Z0 => UQVN_N205, A0 => A13, A1 => UQVN_N224, A2 => B14);
UQVB_B254 : AND4
	PORT MAP (Z0 => UQVN_N204, A0 => B12, A1 => B13, A2 => UQVN_N225, 
	A3 => UQVN_N238);
UQVB_B255 : OR12
	PORT MAP (Z0 => UQVN_N219, A0 => UQVN_N215, A1 => UQVN_N214, A2 => UQVN_N213, 
	A3 => UQVN_N212, A4 => UQVN_N211, A5 => UQVN_N210, A6 => UQVN_N209, 
	A7 => UQVN_N208, A8 => UQVN_N207, A9 => UQVN_N206, A10 => UQVN_N205, 
	A11 => UQVN_N204);
UQVB_B256 : OR3
	PORT MAP (Z0 => UQVN_N217, A0 => UQVN_N216, A1 => UQVN_N218, A2 => UQVN_N219);
UQVB_B257 : XOR2
	PORT MAP (Z0 => Z15, A0 => A15, A1 => UQVN_N230);
UQVB_B258 : AND2
	PORT MAP (Z0 => UQVN_N229, A0 => UQVN_N235, A1 => UQVN_N239);
UQVB_B259 : AND2
	PORT MAP (Z0 => UQVN_N228, A0 => B15, A1 => UQVN_N227);
UQVB_B260 : OR2
	PORT MAP (Z0 => UQVN_N230, A0 => UQVN_N228, A1 => UQVN_N229);
UQVB_B261 : INV
	PORT MAP (ZN0 => UQVN_N231, A0 => A15);
UQVB_B262 : INV
	PORT MAP (ZN0 => UQVN_N235, A0 => B15);
UQVB_B263 : INV
	PORT MAP (ZN0 => UQVN_N227, A0 => UQVN_N239);
UQVB_B264 : AND2
	PORT MAP (Z0 => UQVN_N232, A0 => UQVN_N239, A1 => B15);
UQVB_B265 : AND2
	PORT MAP (Z0 => UQVN_N233, A0 => UQVN_N239, A1 => UQVN_N231);
UQVB_B266 : AND2
	PORT MAP (Z0 => UQVN_N234, A0 => B15, A1 => UQVN_N231);
UQVB_B267 : OR3
	PORT MAP (Z0 => BO, A0 => UQVN_N232, A1 => UQVN_N233, A2 => UQVN_N234);
END lattice_arch;
-- VHDL netlist for SUBF2
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBF2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        BI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBF2;


ARCHITECTURE lattice_arch OF SUBF2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => BI);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => BI, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => BI, A1 => UQVN_N19, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => BI, A1 => UQVN_N18, A2 => B1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => BI, A1 => B1, A2 => B0);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N19, A1 => UQVN_N18, A2 => B0);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N18, A1 => B1, A2 => B0);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N19, A1 => B1);
UQVB_B9 : OR7
	PORT MAP (Z0 => BO, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N5, A5 => UQVN_N7, A6 => UQVN_N6);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => B1, A2 => UQVN_N22);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B1, A1 => UQVN_N20, A2 => UQVN_N22);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N18, A1 => UQVN_N21, A2 => BI);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N21, A1 => B0, A2 => BI);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => A0, A1 => B1, A2 => UQVN_N20);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N18, A1 => UQVN_N21, A2 => B0);
UQVB_B16 : OR6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N12, A5 => UQVN_N13);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N14);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => B0);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => B1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => A1);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => A0);
UQVB_B22 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N15);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N16, A1 => UQVN_N17);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => BI);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N22, A1 => B0);
END lattice_arch;
-- VHDL netlist for SUBF4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBF4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        BI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBF4;


ARCHITECTURE lattice_arch OF SUBF4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => BI);
UQVB_B2 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => BI, A1 => UQVN_N19, A2 => UQVN_N18);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N2, A0 => BI, A1 => UQVN_N19, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N1, A0 => BI, A1 => UQVN_N18, A2 => B1);
UQVB_B5 : AND3
	PORT MAP (Z0 => UQVN_N4, A0 => BI, A1 => B1, A2 => B0);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N19, A1 => UQVN_N18, A2 => B0);
UQVB_B7 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N18, A1 => B1, A2 => B0);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N19, A1 => B1);
UQVB_B9 : OR7
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N3, A1 => UQVN_N2, A2 => UQVN_N1, 
	A3 => UQVN_N4, A4 => UQVN_N5, A5 => UQVN_N7, A6 => UQVN_N6);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A0, A1 => B1, A2 => UQVN_N22);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B1, A1 => UQVN_N20, A2 => UQVN_N22);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N18, A1 => UQVN_N21, A2 => BI);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N21, A1 => B0, A2 => BI);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => A0, A1 => B1, A2 => UQVN_N20);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N18, A1 => UQVN_N21, A2 => B0);
UQVB_B16 : OR6
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N8, A1 => UQVN_N9, A2 => UQVN_N10, 
	A3 => UQVN_N11, A4 => UQVN_N12, A5 => UQVN_N13);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N14);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N20, A0 => B0);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => B1);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N19, A0 => A1);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => A0);
UQVB_B22 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N15);
UQVB_B23 : OR2
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N16, A1 => UQVN_N17);
UQVB_B24 : AND2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => BI);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N22, A1 => B0);
UQVB_B26 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => UQVN_N45);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N45, A1 => UQVN_N41, A2 => UQVN_N40);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N45, A1 => UQVN_N41, A2 => B2);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N45, A1 => UQVN_N40, A2 => B3);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N45, A1 => B3, A2 => B2);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N41, A1 => UQVN_N40, A2 => B2);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N40, A1 => B3, A2 => B2);
UQVB_B33 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N41, A1 => B3);
UQVB_B34 : OR7
	PORT MAP (Z0 => BO, A0 => UQVN_N25, A1 => UQVN_N24, A2 => UQVN_N23, 
	A3 => UQVN_N26, A4 => UQVN_N27, A5 => UQVN_N29, A6 => UQVN_N28);
UQVB_B35 : AND3
	PORT MAP (Z0 => UQVN_N30, A0 => A2, A1 => B3, A2 => UQVN_N44);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N31, A0 => B3, A1 => UQVN_N42, A2 => UQVN_N44);
UQVB_B37 : AND3
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N40, A1 => UQVN_N43, A2 => UQVN_N45);
UQVB_B38 : AND3
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N43, A1 => B2, A2 => UQVN_N45);
UQVB_B39 : AND3
	PORT MAP (Z0 => UQVN_N34, A0 => A2, A1 => B3, A2 => UQVN_N42);
UQVB_B40 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N40, A1 => UQVN_N43, A2 => B2);
UQVB_B41 : OR6
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N30, A1 => UQVN_N31, A2 => UQVN_N32, 
	A3 => UQVN_N33, A4 => UQVN_N34, A5 => UQVN_N35);
UQVB_B42 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N36);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B2);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => B3);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => A3);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => A2);
UQVB_B47 : XOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N37);
UQVB_B48 : OR2
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N38, A1 => UQVN_N39);
UQVB_B49 : AND2
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N42, A1 => UQVN_N45);
UQVB_B50 : AND2
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N44, A1 => B2);
END lattice_arch;
-- VHDL netlist for SUBF8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBF8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        BI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBF8;


ARCHITECTURE lattice_arch OF SUBF8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 G0, G1, G2, G3,
	 G4, G5, G6, G7,
	 P0, P1, P2, P3,
	 P4, P5, P6, P7 : std_logic;


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


BEGIN

UQVB_B1 : XOR2
	PORT MAP (Z0 => P7, A0 => A7, A1 => B7);
UQVB_B2 : XOR2
	PORT MAP (Z0 => P6, A0 => A6, A1 => B6);
UQVB_B3 : XOR2
	PORT MAP (Z0 => P5, A0 => A5, A1 => B5);
UQVB_B4 : XOR2
	PORT MAP (Z0 => P4, A0 => A4, A1 => B4);
UQVB_B5 : XOR2
	PORT MAP (Z0 => P3, A0 => A3, A1 => B3);
UQVB_B6 : XOR2
	PORT MAP (Z0 => P2, A0 => A2, A1 => B2);
UQVB_B7 : XOR2
	PORT MAP (Z0 => P1, A0 => A1, A1 => B1);
UQVB_B8 : XOR2
	PORT MAP (Z0 => P0, A0 => A0, A1 => B0);
UQVB_B9 : AND2
	PORT MAP (Z0 => G7, A0 => UQVN_N8, A1 => B7);
UQVB_B10 : AND2
	PORT MAP (Z0 => G6, A0 => UQVN_N7, A1 => B6);
UQVB_B11 : AND2
	PORT MAP (Z0 => G5, A0 => UQVN_N6, A1 => B5);
UQVB_B12 : AND2
	PORT MAP (Z0 => G4, A0 => UQVN_N5, A1 => B4);
UQVB_B13 : AND2
	PORT MAP (Z0 => G3, A0 => UQVN_N4, A1 => B3);
UQVB_B14 : AND2
	PORT MAP (Z0 => G2, A0 => UQVN_N3, A1 => B2);
UQVB_B15 : AND2
	PORT MAP (Z0 => G1, A0 => UQVN_N2, A1 => B1);
UQVB_B16 : AND2
	PORT MAP (Z0 => G0, A0 => UQVN_N1, A1 => B0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N1, A0 => A0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => A1);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => A2);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => A3);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => A4);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => A5);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => A6);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => A7);
UQVB_B25 : AND8
	PORT MAP (Z0 => UQVN_N32, A0 => G0, A1 => UQVN_N30, A2 => UQVN_N29, 
	A3 => UQVN_N28, A4 => UQVN_N27, A5 => UQVN_N26, A6 => UQVN_N25, 
	A7 => UQVN_N22);
UQVB_B26 : OR6
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N13, A1 => UQVN_N12, A2 => UQVN_N11, 
	A3 => UQVN_N14, A4 => UQVN_N15, A5 => G4);
UQVB_B27 : LXOR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N16, A1 => P5);
UQVB_B28 : AND7
	PORT MAP (Z0 => UQVN_N31, A0 => G1, A1 => UQVN_N29, A2 => UQVN_N28, 
	A3 => UQVN_N27, A4 => UQVN_N26, A5 => UQVN_N25, A6 => UQVN_N22);
UQVB_B29 : OR5
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N36, A1 => UQVN_N35, A2 => UQVN_N38, 
	A3 => UQVN_N37, A4 => G7);
UQVB_B30 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => G0, A1 => UQVN_N17);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => BI, A1 => UQVN_N18, A2 => UQVN_N17);
UQVB_B32 : OR3
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N19, A1 => UQVN_N20, A2 => G1);
UQVB_B33 : AND9
	PORT MAP (Z0 => UQVN_N34, A0 => BI, A1 => UQVN_N23, A2 => UQVN_N30, 
	A3 => UQVN_N29, A4 => UQVN_N28, A5 => UQVN_N27, A6 => UQVN_N26, 
	A7 => UQVN_N25, A8 => UQVN_N22);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N21, A1 => P2);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => P7);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => P6);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => P5);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => P4);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => P3);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => P2);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => P1);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => P0);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => P0);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => P1);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => P2);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => P3);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => P4);
UQVB_B48 : AND6
	PORT MAP (Z0 => UQVN_N33, A0 => G2, A1 => UQVN_N28, A2 => UQVN_N27, 
	A3 => UQVN_N26, A4 => UQVN_N25, A5 => UQVN_N22);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => P1);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N18, A0 => P0);
UQVB_B51 : AND5
	PORT MAP (Z0 => UQVN_N36, A0 => G3, A1 => UQVN_N27, A2 => UQVN_N26, 
	A3 => UQVN_N25, A4 => UQVN_N22);
UQVB_B52 : AND2
	PORT MAP (Z0 => UQVN_N37, A0 => G6, A1 => UQVN_N22);
UQVB_B53 : AND3
	PORT MAP (Z0 => UQVN_N38, A0 => G5, A1 => UQVN_N25, A2 => UQVN_N22);
UQVB_B54 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => G4, A1 => UQVN_N26, A2 => UQVN_N25, 
	A3 => UQVN_N22);
UQVB_B55 : OR4
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N34, A1 => UQVN_N32, A2 => UQVN_N31, 
	A3 => UQVN_N33);
UQVB_B56 : OR2
	PORT MAP (Z0 => BO, A0 => UQVN_N40, A1 => UQVN_N39);
UQVB_B57 : AND6
	PORT MAP (Z0 => UQVN_N13, A0 => BI, A1 => UQVN_N24, A2 => UQVN_N10, 
	A3 => UQVN_N9, A4 => UQVN_N42, A5 => UQVN_N41);
UQVB_B58 : AND5
	PORT MAP (Z0 => UQVN_N12, A0 => G0, A1 => UQVN_N10, A2 => UQVN_N9, 
	A3 => UQVN_N42, A4 => UQVN_N41);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => G1, A1 => UQVN_N9, A2 => UQVN_N42, 
	A3 => UQVN_N41);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => G2, A1 => UQVN_N42, A2 => UQVN_N41);
UQVB_B61 : AND2
	PORT MAP (Z0 => UQVN_N15, A0 => G3, A1 => UQVN_N41);
UQVB_B62 : AND2
	PORT MAP (Z0 => UQVN_N61, A0 => BI, A1 => UQVN_N43);
UQVB_B63 : OR2
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N61, A1 => G0);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => P6);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => P5);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => P4);
UQVB_B67 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => P3);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => P2);
UQVB_B69 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => P1);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => P0);
UQVB_B71 : OR2
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N51, A1 => UQVN_N50);
UQVB_B72 : LXOR2
	PORT MAP (Z0 => Z1, A0 => UQVN_N60, A1 => P1);
UQVB_B73 : XOR2
	PORT MAP (Z0 => Z0, A0 => BI, A1 => P0);
UQVB_B74 : AND2
	PORT MAP (Z0 => UQVN_N58, A0 => G5, A1 => UQVN_N49);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N56, A0 => G4, A1 => UQVN_N48, A2 => UQVN_N49);
UQVB_B76 : AND4
	PORT MAP (Z0 => UQVN_N57, A0 => G3, A1 => UQVN_N47, A2 => UQVN_N48, 
	A3 => UQVN_N49);
UQVB_B77 : AND5
	PORT MAP (Z0 => UQVN_N54, A0 => G2, A1 => UQVN_N46, A2 => UQVN_N47, 
	A3 => UQVN_N48, A4 => UQVN_N49);
UQVB_B78 : AND6
	PORT MAP (Z0 => UQVN_N52, A0 => G1, A1 => UQVN_N45, A2 => UQVN_N46, 
	A3 => UQVN_N47, A4 => UQVN_N48, A5 => UQVN_N49);
UQVB_B79 : AND7
	PORT MAP (Z0 => UQVN_N53, A0 => G0, A1 => UQVN_N44, A2 => UQVN_N45, 
	A3 => UQVN_N46, A4 => UQVN_N47, A5 => UQVN_N48, A6 => UQVN_N49);
UQVB_B80 : AND8
	PORT MAP (Z0 => UQVN_N55, A0 => BI, A1 => UQVN_N43, A2 => UQVN_N44, 
	A3 => UQVN_N45, A4 => UQVN_N46, A5 => UQVN_N47, A6 => UQVN_N48, 
	A7 => UQVN_N49);
UQVB_B81 : OR5
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N55, A1 => UQVN_N53, A2 => UQVN_N52, 
	A3 => UQVN_N54, A4 => UQVN_N57);
UQVB_B82 : OR3
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N56, A1 => UQVN_N58, A2 => G6);
UQVB_B83 : LXOR2
	PORT MAP (Z0 => Z7, A0 => UQVN_N59, A1 => P7);
UQVB_B84 : AND2
	PORT MAP (Z0 => UQVN_N87, A0 => G2, A1 => UQVN_N90);
UQVB_B85 : AND3
	PORT MAP (Z0 => UQVN_N86, A0 => G1, A1 => UQVN_N91, A2 => UQVN_N90);
UQVB_B86 : AND4
	PORT MAP (Z0 => UQVN_N88, A0 => G0, A1 => UQVN_N62, A2 => UQVN_N91, 
	A3 => UQVN_N90);
UQVB_B87 : AND5
	PORT MAP (Z0 => UQVN_N89, A0 => BI, A1 => UQVN_N71, A2 => UQVN_N62, 
	A3 => UQVN_N91, A4 => UQVN_N90);
UQVB_B88 : OR5
	PORT MAP (Z0 => UQVN_N85, A0 => UQVN_N89, A1 => UQVN_N88, A2 => UQVN_N86, 
	A3 => UQVN_N87, A4 => G3);
UQVB_B89 : LXOR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N63, A1 => P3);
UQVB_B90 : AND2
	PORT MAP (Z0 => UQVN_N68, A0 => G1, A1 => UQVN_N67);
UQVB_B91 : AND3
	PORT MAP (Z0 => UQVN_N65, A0 => G0, A1 => UQVN_N66, A2 => UQVN_N67);
UQVB_B92 : AND4
	PORT MAP (Z0 => UQVN_N64, A0 => BI, A1 => UQVN_N72, A2 => UQVN_N66, 
	A3 => UQVN_N67);
UQVB_B93 : OR4
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N64, A1 => UQVN_N65, A2 => UQVN_N68, 
	A3 => G2);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N76, A0 => P5);
UQVB_B95 : INV
	PORT MAP (ZN0 => UQVN_N75, A0 => P4);
UQVB_B96 : INV
	PORT MAP (ZN0 => UQVN_N74, A0 => P3);
UQVB_B97 : INV
	PORT MAP (ZN0 => UQVN_N73, A0 => P2);
UQVB_B98 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => P1);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => P0);
UQVB_B100 : INV
	PORT MAP (ZN0 => UQVN_N90, A0 => P3);
UQVB_B101 : INV
	PORT MAP (ZN0 => UQVN_N91, A0 => P2);
UQVB_B102 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => P1);
UQVB_B103 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => P0);
UQVB_B104 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => P2);
UQVB_B105 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => P1);
UQVB_B106 : INV
	PORT MAP (ZN0 => UQVN_N72, A0 => P0);
UQVB_B107 : OR2
	PORT MAP (Z0 => UQVN_N92, A0 => UQVN_N78, A1 => UQVN_N77);
UQVB_B108 : OR4
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N82, A1 => UQVN_N80, A2 => UQVN_N79, 
	A3 => UQVN_N81);
UQVB_B109 : LXOR2
	PORT MAP (Z0 => Z4, A0 => UQVN_N85, A1 => P4);
UQVB_B110 : AND2
	PORT MAP (Z0 => UQVN_N83, A0 => G4, A1 => UQVN_N76);
UQVB_B111 : AND3
	PORT MAP (Z0 => UQVN_N84, A0 => G3, A1 => UQVN_N75, A2 => UQVN_N76);
UQVB_B112 : AND4
	PORT MAP (Z0 => UQVN_N81, A0 => G2, A1 => UQVN_N74, A2 => UQVN_N75, 
	A3 => UQVN_N76);
UQVB_B113 : AND5
	PORT MAP (Z0 => UQVN_N79, A0 => G1, A1 => UQVN_N73, A2 => UQVN_N74, 
	A3 => UQVN_N75, A4 => UQVN_N76);
UQVB_B114 : AND6
	PORT MAP (Z0 => UQVN_N80, A0 => G0, A1 => UQVN_N70, A2 => UQVN_N73, 
	A3 => UQVN_N74, A4 => UQVN_N75, A5 => UQVN_N76);
UQVB_B115 : AND7
	PORT MAP (Z0 => UQVN_N82, A0 => BI, A1 => UQVN_N69, A2 => UQVN_N70, 
	A3 => UQVN_N73, A4 => UQVN_N74, A5 => UQVN_N75, A6 => UQVN_N76);
UQVB_B116 : OR3
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N84, A1 => UQVN_N83, A2 => G5);
UQVB_B117 : LXOR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N92, A1 => P6);
END lattice_arch;
-- VHDL netlist for SUBF8A
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBF8A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        BI : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBF8A;


ARCHITECTURE lattice_arch OF SUBF8A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 UQVN_N113, G012, G345, P012,
	 P345 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => P012, A1 => BI);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N112, A0 => G012, A1 => UQVN_N1);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N113, A0 => G345, A1 => UQVN_N2, A2 => UQVN_N3);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => P345, A1 => P012, A2 => BI);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => P345, A1 => G012);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => BI);
UQVB_B7 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => B1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => B2);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => A0);
UQVB_B10 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N43, A1 => BI);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => B0, A1 => UQVN_N46);
UQVB_B12 : OR2
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N4, A1 => UQVN_N5);
UQVB_B13 : LXOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => UQVN_N6);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => A0, A1 => B1, A2 => UQVN_N43);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N44, A1 => B0, A2 => BI);
UQVB_B16 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N40, A1 => UQVN_N44, A2 => BI);
UQVB_B17 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => B1, A1 => UQVN_N43, A2 => UQVN_N46);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => A0, A1 => B1, A2 => UQVN_N46);
UQVB_B19 : OR6
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N10, A1 => UQVN_N9, A2 => UQVN_N7, 
	A3 => UQVN_N8, A4 => UQVN_N12, A5 => UQVN_N11);
UQVB_B20 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N13);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N40, A1 => UQVN_N44, A2 => B0);
UQVB_B22 : AND4
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N40, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N41, A1 => B1, A2 => B2);
UQVB_B24 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N40, A1 => UQVN_N42, A2 => B0, 
	A3 => B1);
UQVB_B25 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N42, A1 => B2);
UQVB_B26 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B0, 
	A3 => B2);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N41, A1 => UQVN_N42, A2 => B1);
UQVB_B28 : AND4
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N40, A1 => UQVN_N41, A2 => UQVN_N42, 
	A3 => B0);
UQVB_B29 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N15, 
	A3 => UQVN_N14, A4 => UQVN_N18, A5 => UQVN_N19, A6 => UQVN_N20);
UQVB_B30 : AND2
	PORT MAP (Z0 => UQVN_N23, A0 => A0, A1 => UQVN_N43);
UQVB_B31 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => A1, A1 => UQVN_N44);
UQVB_B32 : AND2
	PORT MAP (Z0 => UQVN_N22, A0 => A2, A1 => UQVN_N45);
UQVB_B33 : NOR3
	PORT MAP (ZN0 => P012, A0 => UQVN_N23, A1 => UQVN_N21, A2 => UQVN_N22);
UQVB_B34 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => B0);
UQVB_B35 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => A1);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => A2);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N37);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N36, A0 => A0, A1 => A1, A2 => B2, 
	A3 => UQVN_N46);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N40, A1 => UQVN_N41, A2 => UQVN_N45, 
	A3 => BI);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N35, A0 => A0, A1 => A1, A2 => UQVN_N43, 
	A3 => B2);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => A1, A1 => UQVN_N43, A2 => B2, 
	A3 => UQVN_N46);
UQVB_B42 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N40, A1 => UQVN_N41, A2 => B0, 
	A3 => UQVN_N45);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N41, A1 => B0, A2 => UQVN_N45, 
	A3 => BI);
UQVB_B44 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => A0, A1 => UQVN_N44, A2 => B2, 
	A3 => UQVN_N46);
UQVB_B45 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => A0, A1 => UQVN_N43, A2 => UQVN_N44, 
	A3 => B2);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N43, A1 => UQVN_N44, A2 => B2, 
	A3 => UQVN_N46);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N41, A1 => UQVN_N45, A2 => B1);
UQVB_B48 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N40, A1 => B1, A2 => UQVN_N45, 
	A3 => BI);
UQVB_B49 : AND4
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N40, A1 => B0, A2 => B1, 
	A3 => UQVN_N45);
UQVB_B50 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => A1, A1 => UQVN_N44, A2 => B2);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => B0, A1 => B1, A2 => UQVN_N45, 
	A3 => BI);
UQVB_B52 : OR12
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N35, A1 => UQVN_N34, A2 => UQVN_N33, 
	A3 => UQVN_N32, A4 => UQVN_N31, A5 => UQVN_N30, A6 => UQVN_N29, 
	A7 => UQVN_N28, A8 => UQVN_N27, A9 => UQVN_N26, A10 => UQVN_N25, 
	A11 => UQVN_N24);
UQVB_B53 : OR3
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N36, A1 => UQVN_N38, A2 => UQVN_N39);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N89, A0 => UQVN_N112);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N87, A0 => B4);
UQVB_B56 : INV
	PORT MAP (ZN0 => UQVN_N88, A0 => B5);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N83, A0 => A3);
UQVB_B58 : AND2
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N86, A1 => UQVN_N112);
UQVB_B59 : AND2
	PORT MAP (Z0 => UQVN_N48, A0 => B3, A1 => UQVN_N89);
UQVB_B60 : OR2
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N47, A1 => UQVN_N48);
UQVB_B61 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N49);
UQVB_B62 : AND3
	PORT MAP (Z0 => UQVN_N55, A0 => A3, A1 => B4, A2 => UQVN_N86);
UQVB_B63 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N87, A1 => B3, A2 => UQVN_N112);
UQVB_B64 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N83, A1 => UQVN_N87, A2 => UQVN_N112);
UQVB_B65 : AND3
	PORT MAP (Z0 => UQVN_N52, A0 => B4, A1 => UQVN_N86, A2 => UQVN_N89);
UQVB_B66 : AND3
	PORT MAP (Z0 => UQVN_N53, A0 => A3, A1 => B4, A2 => UQVN_N89);
UQVB_B67 : OR6
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N53, A1 => UQVN_N52, A2 => UQVN_N50, 
	A3 => UQVN_N51, A4 => UQVN_N55, A5 => UQVN_N54);
UQVB_B68 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N56);
UQVB_B69 : AND3
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N83, A1 => UQVN_N87, A2 => B3);
UQVB_B70 : AND4
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N83, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B71 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N84, A1 => B4, A2 => B5);
UQVB_B72 : AND4
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N83, A1 => UQVN_N85, A2 => B3, 
	A3 => B4);
UQVB_B73 : AND2
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N85, A1 => B5);
UQVB_B74 : AND4
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N83, A1 => UQVN_N84, A2 => B3, 
	A3 => B5);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N84, A1 => UQVN_N85, A2 => B4);
UQVB_B76 : AND4
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N83, A1 => UQVN_N84, A2 => UQVN_N85, 
	A3 => B3);
UQVB_B77 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N60, A1 => UQVN_N59, A2 => UQVN_N58, 
	A3 => UQVN_N57, A4 => UQVN_N61, A5 => UQVN_N62, A6 => UQVN_N63);
UQVB_B78 : AND2
	PORT MAP (Z0 => UQVN_N66, A0 => A3, A1 => UQVN_N86);
UQVB_B79 : AND2
	PORT MAP (Z0 => UQVN_N64, A0 => A4, A1 => UQVN_N87);
UQVB_B80 : AND2
	PORT MAP (Z0 => UQVN_N65, A0 => A5, A1 => UQVN_N88);
UQVB_B81 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N66, A1 => UQVN_N64, A2 => UQVN_N65);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N86, A0 => B3);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N84, A0 => A4);
UQVB_B84 : INV
	PORT MAP (ZN0 => UQVN_N85, A0 => A5);
UQVB_B85 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N80);
UQVB_B86 : AND4
	PORT MAP (Z0 => UQVN_N79, A0 => A3, A1 => A4, A2 => B5, 
	A3 => UQVN_N89);
UQVB_B87 : AND4
	PORT MAP (Z0 => UQVN_N81, A0 => UQVN_N83, A1 => UQVN_N84, A2 => UQVN_N88, 
	A3 => UQVN_N112);
UQVB_B88 : AND4
	PORT MAP (Z0 => UQVN_N78, A0 => A3, A1 => A4, A2 => UQVN_N86, 
	A3 => B5);
UQVB_B89 : AND4
	PORT MAP (Z0 => UQVN_N77, A0 => A4, A1 => UQVN_N86, A2 => B5, 
	A3 => UQVN_N89);
UQVB_B90 : AND4
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N83, A1 => UQVN_N84, A2 => B3, 
	A3 => UQVN_N88);
UQVB_B91 : AND4
	PORT MAP (Z0 => UQVN_N75, A0 => UQVN_N84, A1 => B3, A2 => UQVN_N88, 
	A3 => UQVN_N112);
UQVB_B92 : AND4
	PORT MAP (Z0 => UQVN_N74, A0 => A3, A1 => UQVN_N87, A2 => B5, 
	A3 => UQVN_N89);
UQVB_B93 : AND4
	PORT MAP (Z0 => UQVN_N73, A0 => A3, A1 => UQVN_N86, A2 => UQVN_N87, 
	A3 => B5);
UQVB_B94 : AND4
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N86, A1 => UQVN_N87, A2 => B5, 
	A3 => UQVN_N89);
UQVB_B95 : AND3
	PORT MAP (Z0 => UQVN_N71, A0 => UQVN_N84, A1 => UQVN_N88, A2 => B4);
UQVB_B96 : AND4
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N83, A1 => B4, A2 => UQVN_N88, 
	A3 => UQVN_N112);
UQVB_B97 : AND4
	PORT MAP (Z0 => UQVN_N69, A0 => UQVN_N83, A1 => B3, A2 => B4, 
	A3 => UQVN_N88);
UQVB_B98 : AND3
	PORT MAP (Z0 => UQVN_N68, A0 => A4, A1 => UQVN_N87, A2 => B5);
UQVB_B99 : AND4
	PORT MAP (Z0 => UQVN_N67, A0 => B3, A1 => B4, A2 => UQVN_N88, 
	A3 => UQVN_N112);
UQVB_B100 : OR12
	PORT MAP (Z0 => UQVN_N82, A0 => UQVN_N78, A1 => UQVN_N77, A2 => UQVN_N76, 
	A3 => UQVN_N75, A4 => UQVN_N74, A5 => UQVN_N73, A6 => UQVN_N72, 
	A7 => UQVN_N71, A8 => UQVN_N70, A9 => UQVN_N69, A10 => UQVN_N68, 
	A11 => UQVN_N67);
UQVB_B101 : OR3
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N79, A1 => UQVN_N81, A2 => UQVN_N82);
UQVB_B102 : INV
	PORT MAP (ZN0 => UQVN_N111, A0 => UQVN_N113);
UQVB_B103 : AND3
	PORT MAP (Z0 => UQVN_N92, A0 => UQVN_N113, A1 => UQVN_N108, A2 => UQVN_N107);
UQVB_B104 : AND3
	PORT MAP (Z0 => UQVN_N91, A0 => UQVN_N113, A1 => UQVN_N108, A2 => B6);
UQVB_B105 : AND3
	PORT MAP (Z0 => UQVN_N90, A0 => UQVN_N113, A1 => UQVN_N107, A2 => B7);
UQVB_B106 : AND3
	PORT MAP (Z0 => UQVN_N93, A0 => UQVN_N113, A1 => B7, A2 => B6);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N94, A0 => UQVN_N108, A1 => UQVN_N107, A2 => B6);
UQVB_B108 : AND3
	PORT MAP (Z0 => UQVN_N96, A0 => UQVN_N107, A1 => B7, A2 => B6);
UQVB_B109 : AND2
	PORT MAP (Z0 => UQVN_N95, A0 => UQVN_N108, A1 => B7);
UQVB_B110 : OR7
	PORT MAP (Z0 => BO, A0 => UQVN_N92, A1 => UQVN_N91, A2 => UQVN_N90, 
	A3 => UQVN_N93, A4 => UQVN_N94, A5 => UQVN_N96, A6 => UQVN_N95);
UQVB_B111 : AND3
	PORT MAP (Z0 => UQVN_N97, A0 => A6, A1 => B7, A2 => UQVN_N111);
UQVB_B112 : AND3
	PORT MAP (Z0 => UQVN_N98, A0 => B7, A1 => UQVN_N109, A2 => UQVN_N111);
UQVB_B113 : AND3
	PORT MAP (Z0 => UQVN_N99, A0 => UQVN_N107, A1 => UQVN_N110, A2 => UQVN_N113);
UQVB_B114 : AND3
	PORT MAP (Z0 => UQVN_N100, A0 => UQVN_N110, A1 => B6, A2 => UQVN_N113);
UQVB_B115 : AND3
	PORT MAP (Z0 => UQVN_N101, A0 => A6, A1 => B7, A2 => UQVN_N109);
UQVB_B116 : AND3
	PORT MAP (Z0 => UQVN_N102, A0 => UQVN_N107, A1 => UQVN_N110, A2 => B6);
UQVB_B117 : OR6
	PORT MAP (Z0 => UQVN_N103, A0 => UQVN_N97, A1 => UQVN_N98, A2 => UQVN_N99, 
	A3 => UQVN_N100, A4 => UQVN_N101, A5 => UQVN_N102);
UQVB_B118 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N103);
UQVB_B119 : INV
	PORT MAP (ZN0 => UQVN_N109, A0 => B6);
UQVB_B120 : INV
	PORT MAP (ZN0 => UQVN_N110, A0 => B7);
UQVB_B121 : INV
	PORT MAP (ZN0 => UQVN_N108, A0 => A7);
UQVB_B122 : INV
	PORT MAP (ZN0 => UQVN_N107, A0 => A6);
UQVB_B123 : XOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N104);
UQVB_B124 : OR2
	PORT MAP (Z0 => UQVN_N104, A0 => UQVN_N105, A1 => UQVN_N106);
UQVB_B125 : AND2
	PORT MAP (Z0 => UQVN_N105, A0 => UQVN_N109, A1 => UQVN_N113);
UQVB_B126 : AND2
	PORT MAP (Z0 => UQVN_N106, A0 => UQVN_N111, A1 => B6);
END lattice_arch;
-- VHDL netlist for SUBH1
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH1 IS 
    PORT (
        A0 : IN std_logic;
        B0 : IN std_logic;
        Z0 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBH1;


ARCHITECTURE lattice_arch OF SUBH1 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N4, A1 => B0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N3, A1 => A0);
UQVB_B3 : AND2
	PORT MAP (Z0 => BO, A0 => B0, A1 => UQVN_N4);
UQVB_B4 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N1, A1 => UQVN_N2);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => B0);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => A0);
END lattice_arch;
-- VHDL netlist for SUBH16A
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH16A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        A12 : IN std_logic;
        A13 : IN std_logic;
        A14 : IN std_logic;
        A15 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B10 : IN std_logic;
        B11 : IN std_logic;
        B12 : IN std_logic;
        B13 : IN std_logic;
        B14 : IN std_logic;
        B15 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        B8 : IN std_logic;
        B9 : IN std_logic;
        BO : OUT std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z10 : OUT std_logic;
        Z11 : OUT std_logic;
        Z12 : OUT std_logic;
        Z13 : OUT std_logic;
        Z14 : OUT std_logic;
        Z15 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        Z8 : OUT std_logic;
        Z9 : OUT std_logic
    );
END SUBH16A;


ARCHITECTURE lattice_arch OF SUBH16A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, UQVN_N94, UQVN_N95, UQVN_N96,
	 UQVN_N97, UQVN_N98, UQVN_N99, UQVN_N100,
	 UQVN_N101, UQVN_N102, UQVN_N103, UQVN_N104,
	 UQVN_N105, UQVN_N106, UQVN_N107, UQVN_N108,
	 UQVN_N109, UQVN_N110, UQVN_N111, UQVN_N112,
	 UQVN_N113, UQVN_N114, UQVN_N115, UQVN_N116,
	 UQVN_N117, UQVN_N118, UQVN_N119, UQVN_N120,
	 UQVN_N121, UQVN_N122, UQVN_N123, UQVN_N124,
	 UQVN_N125, UQVN_N126, UQVN_N127, UQVN_N128,
	 UQVN_N129, UQVN_N130, UQVN_N131, UQVN_N132,
	 UQVN_N133, UQVN_N134, UQVN_N135, UQVN_N136,
	 UQVN_N137, UQVN_N138, UQVN_N139, UQVN_N140,
	 UQVN_N141, UQVN_N142, UQVN_N143, UQVN_N144,
	 UQVN_N145, UQVN_N146, UQVN_N147, UQVN_N148,
	 UQVN_N149, UQVN_N150, UQVN_N151, UQVN_N152,
	 UQVN_N153, UQVN_N154, UQVN_N155, UQVN_N156,
	 UQVN_N157, UQVN_N158, UQVN_N159, UQVN_N160,
	 UQVN_N161, UQVN_N162, UQVN_N163, UQVN_N164,
	 UQVN_N165, UQVN_N166, UQVN_N167, UQVN_N168,
	 UQVN_N169, UQVN_N170, UQVN_N171, UQVN_N172,
	 UQVN_N173, UQVN_N174, UQVN_N175, UQVN_N176,
	 UQVN_N177, UQVN_N178, UQVN_N179, UQVN_N180,
	 UQVN_N181, UQVN_N182, UQVN_N183, UQVN_N184,
	 UQVN_N185, UQVN_N186, UQVN_N187, UQVN_N188,
	 UQVN_N189, UQVN_N190, UQVN_N191, UQVN_N192,
	 UQVN_N193, UQVN_N194, UQVN_N195, UQVN_N196,
	 UQVN_N197, UQVN_N198, UQVN_N199, UQVN_N200,
	 UQVN_N201, UQVN_N202, UQVN_N203, UQVN_N204,
	 UQVN_N205, UQVN_N206, UQVN_N207, UQVN_N208,
	 UQVN_N209, UQVN_N210, UQVN_N211, UQVN_N212,
	 UQVN_N213, UQVN_N214, UQVN_N215, UQVN_N216,
	 UQVN_N217, UQVN_N218, UQVN_N219, UQVN_N220,
	 UQVN_N221, UQVN_N222, G012, G1214,
	 G345, G911, P1214, P345,
	 P678, P911 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => P345, A1 => G012);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N218, A0 => G345, A1 => UQVN_N1);
UQVB_B3 : OR3
	PORT MAP (Z0 => UQVN_N219, A0 => UQVN_N222, A1 => UQVN_N2, A2 => UQVN_N3);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => P678, A1 => P345, A2 => G012);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => P678, A1 => G345);
UQVB_B6 : OR4
	PORT MAP (Z0 => UQVN_N220, A0 => G911, A1 => UQVN_N4, A2 => UQVN_N5, 
	A3 => UQVN_N6);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => P911, A1 => UQVN_N222);
UQVB_B8 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => P911, A1 => P678, A2 => G345);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => P911, A1 => P678, A2 => P345, 
	A3 => G012);
UQVB_B10 : OR5
	PORT MAP (Z0 => UQVN_N221, A0 => G1214, A1 => UQVN_N7, A2 => UQVN_N8, 
	A3 => UQVN_N9, A4 => UQVN_N10);
UQVB_B11 : AND2
	PORT MAP (Z0 => UQVN_N7, A0 => P1214, A1 => G911);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => P1214, A1 => P911, A2 => UQVN_N222);
UQVB_B13 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => G345);
UQVB_B14 : AND5
	PORT MAP (Z0 => UQVN_N10, A0 => P1214, A1 => P911, A2 => P678, 
	A3 => P345, A4 => G012);
UQVB_B15 : INV
	PORT MAP (ZN0 => UQVN_N53, A0 => G012);
UQVB_B16 : INV
	PORT MAP (ZN0 => UQVN_N51, A0 => B4);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N52, A0 => B5);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N47, A0 => A3);
UQVB_B19 : AND2
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N50, A1 => G012);
UQVB_B20 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => B3, A1 => UQVN_N53);
UQVB_B21 : OR2
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N11, A1 => UQVN_N12);
UQVB_B22 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N13);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => A3, A1 => B4, A2 => UQVN_N50);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N51, A1 => B3, A2 => G012);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N47, A1 => UQVN_N51, A2 => G012);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => B4, A1 => UQVN_N50, A2 => UQVN_N53);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => A3, A1 => B4, A2 => UQVN_N53);
UQVB_B28 : OR6
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N17, A1 => UQVN_N16, A2 => UQVN_N14, 
	A3 => UQVN_N15, A4 => UQVN_N19, A5 => UQVN_N18);
UQVB_B29 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N20);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N47, A1 => UQVN_N51, A2 => B3);
UQVB_B31 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N47, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => UQVN_N48, A1 => B4, A2 => B5);
UQVB_B33 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N47, A1 => UQVN_N49, A2 => B3, 
	A3 => B4);
UQVB_B34 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N49, A1 => B5);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N47, A1 => UQVN_N48, A2 => B3, 
	A3 => B5);
UQVB_B36 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N48, A1 => UQVN_N49, A2 => B4);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N49, 
	A3 => B3);
UQVB_B38 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N24, A1 => UQVN_N23, A2 => UQVN_N22, 
	A3 => UQVN_N21, A4 => UQVN_N25, A5 => UQVN_N26, A6 => UQVN_N27);
UQVB_B39 : AND2
	PORT MAP (Z0 => UQVN_N30, A0 => A3, A1 => UQVN_N50);
UQVB_B40 : AND2
	PORT MAP (Z0 => UQVN_N28, A0 => A4, A1 => UQVN_N51);
UQVB_B41 : AND2
	PORT MAP (Z0 => UQVN_N29, A0 => A5, A1 => UQVN_N52);
UQVB_B42 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N30, A1 => UQVN_N28, A2 => UQVN_N29);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N50, A0 => B3);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N48, A0 => A4);
UQVB_B45 : INV
	PORT MAP (ZN0 => UQVN_N49, A0 => A5);
UQVB_B46 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N44);
UQVB_B47 : AND4
	PORT MAP (Z0 => UQVN_N43, A0 => A3, A1 => A4, A2 => B5, 
	A3 => UQVN_N53);
UQVB_B48 : AND4
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N47, A1 => UQVN_N48, A2 => UQVN_N52, 
	A3 => G012);
UQVB_B49 : AND4
	PORT MAP (Z0 => UQVN_N42, A0 => A3, A1 => A4, A2 => UQVN_N50, 
	A3 => B5);
UQVB_B50 : AND4
	PORT MAP (Z0 => UQVN_N41, A0 => A4, A1 => UQVN_N50, A2 => B5, 
	A3 => UQVN_N53);
UQVB_B51 : AND4
	PORT MAP (Z0 => UQVN_N40, A0 => UQVN_N47, A1 => UQVN_N48, A2 => B3, 
	A3 => UQVN_N52);
UQVB_B52 : AND4
	PORT MAP (Z0 => UQVN_N39, A0 => UQVN_N48, A1 => B3, A2 => UQVN_N52, 
	A3 => G012);
UQVB_B53 : AND4
	PORT MAP (Z0 => UQVN_N38, A0 => A3, A1 => UQVN_N51, A2 => B5, 
	A3 => UQVN_N53);
UQVB_B54 : AND4
	PORT MAP (Z0 => UQVN_N37, A0 => A3, A1 => UQVN_N50, A2 => UQVN_N51, 
	A3 => B5);
UQVB_B55 : AND4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N50, A1 => UQVN_N51, A2 => B5, 
	A3 => UQVN_N53);
UQVB_B56 : AND3
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N48, A1 => UQVN_N52, A2 => B4);
UQVB_B57 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => UQVN_N47, A1 => B4, A2 => UQVN_N52, 
	A3 => G012);
UQVB_B58 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => UQVN_N47, A1 => B3, A2 => B4, 
	A3 => UQVN_N52);
UQVB_B59 : AND3
	PORT MAP (Z0 => UQVN_N32, A0 => A4, A1 => UQVN_N51, A2 => B5);
UQVB_B60 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => B3, A1 => B4, A2 => UQVN_N52, 
	A3 => G012);
UQVB_B61 : OR12
	PORT MAP (Z0 => UQVN_N46, A0 => UQVN_N42, A1 => UQVN_N41, A2 => UQVN_N40, 
	A3 => UQVN_N39, A4 => UQVN_N38, A5 => UQVN_N37, A6 => UQVN_N36, 
	A7 => UQVN_N35, A8 => UQVN_N34, A9 => UQVN_N33, A10 => UQVN_N32, 
	A11 => UQVN_N31);
UQVB_B62 : OR3
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N43, A1 => UQVN_N45, A2 => UQVN_N46);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N96, A0 => UQVN_N218);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N94, A0 => B7);
UQVB_B65 : INV
	PORT MAP (ZN0 => UQVN_N95, A0 => B8);
UQVB_B66 : INV
	PORT MAP (ZN0 => UQVN_N90, A0 => A6);
UQVB_B67 : AND2
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N93, A1 => UQVN_N218);
UQVB_B68 : AND2
	PORT MAP (Z0 => UQVN_N55, A0 => B6, A1 => UQVN_N96);
UQVB_B69 : OR2
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N54, A1 => UQVN_N55);
UQVB_B70 : LXOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N56);
UQVB_B71 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => A6, A1 => B7, A2 => UQVN_N93);
UQVB_B72 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N94, A1 => B6, A2 => UQVN_N218);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N90, A1 => UQVN_N94, A2 => UQVN_N218);
UQVB_B74 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => B7, A1 => UQVN_N93, A2 => UQVN_N96);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N60, A0 => A6, A1 => B7, A2 => UQVN_N96);
UQVB_B76 : OR6
	PORT MAP (Z0 => UQVN_N63, A0 => UQVN_N60, A1 => UQVN_N59, A2 => UQVN_N57, 
	A3 => UQVN_N58, A4 => UQVN_N62, A5 => UQVN_N61);
UQVB_B77 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N63);
UQVB_B78 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N90, A1 => UQVN_N94, A2 => B6);
UQVB_B79 : AND4
	PORT MAP (Z0 => UQVN_N67, A0 => UQVN_N90, A1 => B6, A2 => B7, 
	A3 => B8);
UQVB_B80 : AND3
	PORT MAP (Z0 => UQVN_N66, A0 => UQVN_N91, A1 => B7, A2 => B8);
UQVB_B81 : AND4
	PORT MAP (Z0 => UQVN_N65, A0 => UQVN_N90, A1 => UQVN_N92, A2 => B6, 
	A3 => B7);
UQVB_B82 : AND2
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N92, A1 => B8);
UQVB_B83 : AND4
	PORT MAP (Z0 => UQVN_N68, A0 => UQVN_N90, A1 => UQVN_N91, A2 => B6, 
	A3 => B8);
UQVB_B84 : AND3
	PORT MAP (Z0 => UQVN_N69, A0 => UQVN_N91, A1 => UQVN_N92, A2 => B7);
UQVB_B85 : AND4
	PORT MAP (Z0 => UQVN_N70, A0 => UQVN_N90, A1 => UQVN_N91, A2 => UQVN_N92, 
	A3 => B6);
UQVB_B86 : OR7
	PORT MAP (Z0 => UQVN_N222, A0 => UQVN_N67, A1 => UQVN_N66, A2 => UQVN_N65, 
	A3 => UQVN_N64, A4 => UQVN_N68, A5 => UQVN_N69, A6 => UQVN_N70);
UQVB_B87 : AND2
	PORT MAP (Z0 => UQVN_N73, A0 => A6, A1 => UQVN_N93);
UQVB_B88 : AND2
	PORT MAP (Z0 => UQVN_N71, A0 => A7, A1 => UQVN_N94);
UQVB_B89 : AND2
	PORT MAP (Z0 => UQVN_N72, A0 => A8, A1 => UQVN_N95);
UQVB_B90 : NOR3
	PORT MAP (ZN0 => P678, A0 => UQVN_N73, A1 => UQVN_N71, A2 => UQVN_N72);
UQVB_B91 : INV
	PORT MAP (ZN0 => UQVN_N93, A0 => B6);
UQVB_B92 : INV
	PORT MAP (ZN0 => UQVN_N91, A0 => A7);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N92, A0 => A8);
UQVB_B94 : LXOR2
	PORT MAP (Z0 => Z8, A0 => A8, A1 => UQVN_N87);
UQVB_B95 : AND4
	PORT MAP (Z0 => UQVN_N86, A0 => A6, A1 => A7, A2 => B8, 
	A3 => UQVN_N96);
UQVB_B96 : AND4
	PORT MAP (Z0 => UQVN_N88, A0 => UQVN_N90, A1 => UQVN_N91, A2 => UQVN_N95, 
	A3 => UQVN_N218);
UQVB_B97 : AND4
	PORT MAP (Z0 => UQVN_N85, A0 => A6, A1 => A7, A2 => UQVN_N93, 
	A3 => B8);
UQVB_B98 : AND4
	PORT MAP (Z0 => UQVN_N84, A0 => A7, A1 => UQVN_N93, A2 => B8, 
	A3 => UQVN_N96);
UQVB_B99 : AND4
	PORT MAP (Z0 => UQVN_N83, A0 => UQVN_N90, A1 => UQVN_N91, A2 => B6, 
	A3 => UQVN_N95);
UQVB_B100 : AND4
	PORT MAP (Z0 => UQVN_N82, A0 => UQVN_N91, A1 => B6, A2 => UQVN_N95, 
	A3 => UQVN_N218);
UQVB_B101 : AND4
	PORT MAP (Z0 => UQVN_N81, A0 => A6, A1 => UQVN_N94, A2 => B8, 
	A3 => UQVN_N96);
UQVB_B102 : AND4
	PORT MAP (Z0 => UQVN_N80, A0 => A6, A1 => UQVN_N93, A2 => UQVN_N94, 
	A3 => B8);
UQVB_B103 : AND4
	PORT MAP (Z0 => UQVN_N79, A0 => UQVN_N93, A1 => UQVN_N94, A2 => B8, 
	A3 => UQVN_N96);
UQVB_B104 : AND3
	PORT MAP (Z0 => UQVN_N78, A0 => UQVN_N91, A1 => UQVN_N95, A2 => B7);
UQVB_B105 : AND4
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N90, A1 => B7, A2 => UQVN_N95, 
	A3 => UQVN_N218);
UQVB_B106 : AND4
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N90, A1 => B6, A2 => B7, 
	A3 => UQVN_N95);
UQVB_B107 : AND3
	PORT MAP (Z0 => UQVN_N75, A0 => A7, A1 => UQVN_N94, A2 => B8);
UQVB_B108 : AND4
	PORT MAP (Z0 => UQVN_N74, A0 => B6, A1 => B7, A2 => UQVN_N95, 
	A3 => UQVN_N218);
UQVB_B109 : OR12
	PORT MAP (Z0 => UQVN_N89, A0 => UQVN_N85, A1 => UQVN_N84, A2 => UQVN_N83, 
	A3 => UQVN_N82, A4 => UQVN_N81, A5 => UQVN_N80, A6 => UQVN_N79, 
	A7 => UQVN_N78, A8 => UQVN_N77, A9 => UQVN_N76, A10 => UQVN_N75, 
	A11 => UQVN_N74);
UQVB_B110 : OR3
	PORT MAP (Z0 => UQVN_N87, A0 => UQVN_N86, A1 => UQVN_N88, A2 => UQVN_N89);
UQVB_B111 : INV
	PORT MAP (ZN0 => UQVN_N139, A0 => UQVN_N219);
UQVB_B112 : INV
	PORT MAP (ZN0 => UQVN_N137, A0 => B10);
UQVB_B113 : INV
	PORT MAP (ZN0 => UQVN_N138, A0 => B11);
UQVB_B114 : INV
	PORT MAP (ZN0 => UQVN_N133, A0 => A9);
UQVB_B115 : AND2
	PORT MAP (Z0 => UQVN_N97, A0 => UQVN_N136, A1 => UQVN_N219);
UQVB_B116 : AND2
	PORT MAP (Z0 => UQVN_N98, A0 => B9, A1 => UQVN_N139);
UQVB_B117 : OR2
	PORT MAP (Z0 => UQVN_N99, A0 => UQVN_N97, A1 => UQVN_N98);
UQVB_B118 : LXOR2
	PORT MAP (Z0 => Z9, A0 => A9, A1 => UQVN_N99);
UQVB_B119 : AND3
	PORT MAP (Z0 => UQVN_N105, A0 => A9, A1 => B10, A2 => UQVN_N136);
UQVB_B120 : AND3
	PORT MAP (Z0 => UQVN_N101, A0 => UQVN_N137, A1 => B9, A2 => UQVN_N219);
UQVB_B121 : AND3
	PORT MAP (Z0 => UQVN_N100, A0 => UQVN_N133, A1 => UQVN_N137, A2 => UQVN_N219);
UQVB_B122 : AND3
	PORT MAP (Z0 => UQVN_N102, A0 => B10, A1 => UQVN_N136, A2 => UQVN_N139);
UQVB_B123 : AND3
	PORT MAP (Z0 => UQVN_N103, A0 => A9, A1 => B10, A2 => UQVN_N139);
UQVB_B124 : OR6
	PORT MAP (Z0 => UQVN_N106, A0 => UQVN_N103, A1 => UQVN_N102, A2 => UQVN_N100, 
	A3 => UQVN_N101, A4 => UQVN_N105, A5 => UQVN_N104);
UQVB_B125 : LXOR2
	PORT MAP (Z0 => Z10, A0 => A10, A1 => UQVN_N106);
UQVB_B126 : AND3
	PORT MAP (Z0 => UQVN_N104, A0 => UQVN_N133, A1 => UQVN_N137, A2 => B9);
UQVB_B127 : AND4
	PORT MAP (Z0 => UQVN_N110, A0 => UQVN_N133, A1 => B9, A2 => B10, 
	A3 => B11);
UQVB_B128 : AND3
	PORT MAP (Z0 => UQVN_N109, A0 => UQVN_N134, A1 => B10, A2 => B11);
UQVB_B129 : AND4
	PORT MAP (Z0 => UQVN_N108, A0 => UQVN_N133, A1 => UQVN_N135, A2 => B9, 
	A3 => B10);
UQVB_B130 : AND2
	PORT MAP (Z0 => UQVN_N107, A0 => UQVN_N135, A1 => B11);
UQVB_B131 : AND4
	PORT MAP (Z0 => UQVN_N111, A0 => UQVN_N133, A1 => UQVN_N134, A2 => B9, 
	A3 => B11);
UQVB_B132 : AND3
	PORT MAP (Z0 => UQVN_N112, A0 => UQVN_N134, A1 => UQVN_N135, A2 => B10);
UQVB_B133 : AND4
	PORT MAP (Z0 => UQVN_N113, A0 => UQVN_N133, A1 => UQVN_N134, A2 => UQVN_N135, 
	A3 => B9);
UQVB_B134 : OR7
	PORT MAP (Z0 => G911, A0 => UQVN_N110, A1 => UQVN_N109, A2 => UQVN_N108, 
	A3 => UQVN_N107, A4 => UQVN_N111, A5 => UQVN_N112, A6 => UQVN_N113);
UQVB_B135 : AND2
	PORT MAP (Z0 => UQVN_N116, A0 => A9, A1 => UQVN_N136);
UQVB_B136 : AND2
	PORT MAP (Z0 => UQVN_N114, A0 => A10, A1 => UQVN_N137);
UQVB_B137 : AND2
	PORT MAP (Z0 => UQVN_N115, A0 => A11, A1 => UQVN_N138);
UQVB_B138 : NOR3
	PORT MAP (ZN0 => P911, A0 => UQVN_N116, A1 => UQVN_N114, A2 => UQVN_N115);
UQVB_B139 : INV
	PORT MAP (ZN0 => UQVN_N136, A0 => B9);
UQVB_B140 : INV
	PORT MAP (ZN0 => UQVN_N134, A0 => A10);
UQVB_B141 : INV
	PORT MAP (ZN0 => UQVN_N135, A0 => A11);
UQVB_B142 : LXOR2
	PORT MAP (Z0 => Z11, A0 => A11, A1 => UQVN_N130);
UQVB_B143 : AND4
	PORT MAP (Z0 => UQVN_N129, A0 => A9, A1 => A10, A2 => B11, 
	A3 => UQVN_N139);
UQVB_B144 : AND4
	PORT MAP (Z0 => UQVN_N131, A0 => UQVN_N133, A1 => UQVN_N134, A2 => UQVN_N138, 
	A3 => UQVN_N219);
UQVB_B145 : AND4
	PORT MAP (Z0 => UQVN_N128, A0 => A9, A1 => A10, A2 => UQVN_N136, 
	A3 => B11);
UQVB_B146 : AND4
	PORT MAP (Z0 => UQVN_N127, A0 => A10, A1 => UQVN_N136, A2 => B11, 
	A3 => UQVN_N139);
UQVB_B147 : AND4
	PORT MAP (Z0 => UQVN_N126, A0 => UQVN_N133, A1 => UQVN_N134, A2 => B9, 
	A3 => UQVN_N138);
UQVB_B148 : AND4
	PORT MAP (Z0 => UQVN_N125, A0 => UQVN_N134, A1 => B9, A2 => UQVN_N138, 
	A3 => UQVN_N219);
UQVB_B149 : AND4
	PORT MAP (Z0 => UQVN_N124, A0 => A9, A1 => UQVN_N137, A2 => B11, 
	A3 => UQVN_N139);
UQVB_B150 : AND4
	PORT MAP (Z0 => UQVN_N123, A0 => A9, A1 => UQVN_N136, A2 => UQVN_N137, 
	A3 => B11);
UQVB_B151 : AND4
	PORT MAP (Z0 => UQVN_N122, A0 => UQVN_N136, A1 => UQVN_N137, A2 => B11, 
	A3 => UQVN_N139);
UQVB_B152 : AND3
	PORT MAP (Z0 => UQVN_N121, A0 => UQVN_N134, A1 => UQVN_N138, A2 => B10);
UQVB_B153 : AND4
	PORT MAP (Z0 => UQVN_N120, A0 => UQVN_N133, A1 => B10, A2 => UQVN_N138, 
	A3 => UQVN_N219);
UQVB_B154 : AND4
	PORT MAP (Z0 => UQVN_N119, A0 => UQVN_N133, A1 => B9, A2 => B10, 
	A3 => UQVN_N138);
UQVB_B155 : AND3
	PORT MAP (Z0 => UQVN_N118, A0 => A10, A1 => UQVN_N137, A2 => B11);
UQVB_B156 : AND4
	PORT MAP (Z0 => UQVN_N117, A0 => B9, A1 => B10, A2 => UQVN_N138, 
	A3 => UQVN_N219);
UQVB_B157 : OR12
	PORT MAP (Z0 => UQVN_N132, A0 => UQVN_N128, A1 => UQVN_N127, A2 => UQVN_N126, 
	A3 => UQVN_N125, A4 => UQVN_N124, A5 => UQVN_N123, A6 => UQVN_N122, 
	A7 => UQVN_N121, A8 => UQVN_N120, A9 => UQVN_N119, A10 => UQVN_N118, 
	A11 => UQVN_N117);
UQVB_B158 : OR3
	PORT MAP (Z0 => UQVN_N130, A0 => UQVN_N129, A1 => UQVN_N131, A2 => UQVN_N132);
UQVB_B159 : INV
	PORT MAP (ZN0 => UQVN_N182, A0 => UQVN_N220);
UQVB_B160 : INV
	PORT MAP (ZN0 => UQVN_N180, A0 => B13);
UQVB_B161 : INV
	PORT MAP (ZN0 => UQVN_N181, A0 => B14);
UQVB_B162 : INV
	PORT MAP (ZN0 => UQVN_N176, A0 => A12);
UQVB_B163 : AND2
	PORT MAP (Z0 => UQVN_N140, A0 => UQVN_N179, A1 => UQVN_N220);
UQVB_B164 : AND2
	PORT MAP (Z0 => UQVN_N141, A0 => B12, A1 => UQVN_N182);
UQVB_B165 : OR2
	PORT MAP (Z0 => UQVN_N142, A0 => UQVN_N140, A1 => UQVN_N141);
UQVB_B166 : LXOR2
	PORT MAP (Z0 => Z12, A0 => A12, A1 => UQVN_N142);
UQVB_B167 : AND3
	PORT MAP (Z0 => UQVN_N148, A0 => A12, A1 => B13, A2 => UQVN_N179);
UQVB_B168 : AND3
	PORT MAP (Z0 => UQVN_N144, A0 => UQVN_N180, A1 => B12, A2 => UQVN_N220);
UQVB_B169 : AND3
	PORT MAP (Z0 => UQVN_N143, A0 => UQVN_N176, A1 => UQVN_N180, A2 => UQVN_N220);
UQVB_B170 : AND3
	PORT MAP (Z0 => UQVN_N145, A0 => B13, A1 => UQVN_N179, A2 => UQVN_N182);
UQVB_B171 : AND3
	PORT MAP (Z0 => UQVN_N146, A0 => A12, A1 => B13, A2 => UQVN_N182);
UQVB_B172 : OR6
	PORT MAP (Z0 => UQVN_N149, A0 => UQVN_N146, A1 => UQVN_N145, A2 => UQVN_N143, 
	A3 => UQVN_N144, A4 => UQVN_N148, A5 => UQVN_N147);
UQVB_B173 : LXOR2
	PORT MAP (Z0 => Z13, A0 => A13, A1 => UQVN_N149);
UQVB_B174 : AND3
	PORT MAP (Z0 => UQVN_N147, A0 => UQVN_N176, A1 => UQVN_N180, A2 => B12);
UQVB_B175 : AND4
	PORT MAP (Z0 => UQVN_N153, A0 => UQVN_N176, A1 => B12, A2 => B13, 
	A3 => B14);
UQVB_B176 : AND3
	PORT MAP (Z0 => UQVN_N152, A0 => UQVN_N177, A1 => B13, A2 => B14);
UQVB_B177 : AND4
	PORT MAP (Z0 => UQVN_N151, A0 => UQVN_N176, A1 => UQVN_N178, A2 => B12, 
	A3 => B13);
UQVB_B178 : AND2
	PORT MAP (Z0 => UQVN_N150, A0 => UQVN_N178, A1 => B14);
UQVB_B179 : AND4
	PORT MAP (Z0 => UQVN_N154, A0 => UQVN_N176, A1 => UQVN_N177, A2 => B12, 
	A3 => B14);
UQVB_B180 : AND3
	PORT MAP (Z0 => UQVN_N155, A0 => UQVN_N177, A1 => UQVN_N178, A2 => B13);
UQVB_B181 : AND4
	PORT MAP (Z0 => UQVN_N156, A0 => UQVN_N176, A1 => UQVN_N177, A2 => UQVN_N178, 
	A3 => B12);
UQVB_B182 : OR7
	PORT MAP (Z0 => G1214, A0 => UQVN_N153, A1 => UQVN_N152, A2 => UQVN_N151, 
	A3 => UQVN_N150, A4 => UQVN_N154, A5 => UQVN_N155, A6 => UQVN_N156);
UQVB_B183 : AND2
	PORT MAP (Z0 => UQVN_N159, A0 => A12, A1 => UQVN_N179);
UQVB_B184 : AND2
	PORT MAP (Z0 => UQVN_N157, A0 => A13, A1 => UQVN_N180);
UQVB_B185 : AND2
	PORT MAP (Z0 => UQVN_N158, A0 => A14, A1 => UQVN_N181);
UQVB_B186 : NOR3
	PORT MAP (ZN0 => P1214, A0 => UQVN_N159, A1 => UQVN_N157, A2 => UQVN_N158);
UQVB_B187 : INV
	PORT MAP (ZN0 => UQVN_N179, A0 => B12);
UQVB_B188 : INV
	PORT MAP (ZN0 => UQVN_N177, A0 => A13);
UQVB_B189 : INV
	PORT MAP (ZN0 => UQVN_N178, A0 => A14);
UQVB_B190 : LXOR2
	PORT MAP (Z0 => Z14, A0 => A14, A1 => UQVN_N173);
UQVB_B191 : AND4
	PORT MAP (Z0 => UQVN_N172, A0 => A12, A1 => A13, A2 => B14, 
	A3 => UQVN_N182);
UQVB_B192 : AND4
	PORT MAP (Z0 => UQVN_N174, A0 => UQVN_N176, A1 => UQVN_N177, A2 => UQVN_N181, 
	A3 => UQVN_N220);
UQVB_B193 : AND4
	PORT MAP (Z0 => UQVN_N171, A0 => A12, A1 => A13, A2 => UQVN_N179, 
	A3 => B14);
UQVB_B194 : AND4
	PORT MAP (Z0 => UQVN_N170, A0 => A13, A1 => UQVN_N179, A2 => B14, 
	A3 => UQVN_N182);
UQVB_B195 : AND4
	PORT MAP (Z0 => UQVN_N169, A0 => UQVN_N176, A1 => UQVN_N177, A2 => B12, 
	A3 => UQVN_N181);
UQVB_B196 : AND4
	PORT MAP (Z0 => UQVN_N168, A0 => UQVN_N177, A1 => B12, A2 => UQVN_N181, 
	A3 => UQVN_N220);
UQVB_B197 : AND4
	PORT MAP (Z0 => UQVN_N167, A0 => A12, A1 => UQVN_N180, A2 => B14, 
	A3 => UQVN_N182);
UQVB_B198 : AND4
	PORT MAP (Z0 => UQVN_N166, A0 => A12, A1 => UQVN_N179, A2 => UQVN_N180, 
	A3 => B14);
UQVB_B199 : AND4
	PORT MAP (Z0 => UQVN_N165, A0 => UQVN_N179, A1 => UQVN_N180, A2 => B14, 
	A3 => UQVN_N182);
UQVB_B200 : AND3
	PORT MAP (Z0 => UQVN_N164, A0 => UQVN_N177, A1 => UQVN_N181, A2 => B13);
UQVB_B201 : AND4
	PORT MAP (Z0 => UQVN_N163, A0 => UQVN_N176, A1 => B13, A2 => UQVN_N181, 
	A3 => UQVN_N220);
UQVB_B202 : AND4
	PORT MAP (Z0 => UQVN_N162, A0 => UQVN_N176, A1 => B12, A2 => B13, 
	A3 => UQVN_N181);
UQVB_B203 : AND3
	PORT MAP (Z0 => UQVN_N161, A0 => A13, A1 => UQVN_N180, A2 => B14);
UQVB_B204 : AND4
	PORT MAP (Z0 => UQVN_N160, A0 => B12, A1 => B13, A2 => UQVN_N181, 
	A3 => UQVN_N220);
UQVB_B205 : OR12
	PORT MAP (Z0 => UQVN_N175, A0 => UQVN_N171, A1 => UQVN_N170, A2 => UQVN_N169, 
	A3 => UQVN_N168, A4 => UQVN_N167, A5 => UQVN_N166, A6 => UQVN_N165, 
	A7 => UQVN_N164, A8 => UQVN_N163, A9 => UQVN_N162, A10 => UQVN_N161, 
	A11 => UQVN_N160);
UQVB_B206 : OR3
	PORT MAP (Z0 => UQVN_N173, A0 => UQVN_N172, A1 => UQVN_N174, A2 => UQVN_N175);
UQVB_B207 : INV
	PORT MAP (ZN0 => UQVN_N207, A0 => B1);
UQVB_B208 : INV
	PORT MAP (ZN0 => UQVN_N203, A0 => A0);
UQVB_B209 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N186);
UQVB_B210 : AND3
	PORT MAP (Z0 => UQVN_N185, A0 => UQVN_N203, A1 => B0, A2 => UQVN_N207);
UQVB_B211 : AND4
	PORT MAP (Z0 => UQVN_N190, A0 => UQVN_N203, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B212 : AND3
	PORT MAP (Z0 => UQVN_N189, A0 => UQVN_N204, A1 => B1, A2 => B2);
UQVB_B213 : AND4
	PORT MAP (Z0 => UQVN_N188, A0 => UQVN_N203, A1 => UQVN_N205, A2 => B0, 
	A3 => B1);
UQVB_B214 : AND2
	PORT MAP (Z0 => UQVN_N187, A0 => UQVN_N205, A1 => B2);
UQVB_B215 : AND4
	PORT MAP (Z0 => UQVN_N191, A0 => UQVN_N203, A1 => UQVN_N204, A2 => UQVN_N205, 
	A3 => B0);
UQVB_B216 : AND3
	PORT MAP (Z0 => UQVN_N192, A0 => UQVN_N204, A1 => UQVN_N205, A2 => B1);
UQVB_B217 : AND4
	PORT MAP (Z0 => UQVN_N193, A0 => UQVN_N203, A1 => UQVN_N204, A2 => B0, 
	A3 => B2);
UQVB_B218 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N190, A1 => UQVN_N189, A2 => UQVN_N188, 
	A3 => UQVN_N187, A4 => UQVN_N191, A5 => UQVN_N192, A6 => UQVN_N193);
UQVB_B219 : INV
	PORT MAP (ZN0 => UQVN_N206, A0 => B0);
UQVB_B220 : INV
	PORT MAP (ZN0 => UQVN_N204, A0 => A1);
UQVB_B221 : AND2
	PORT MAP (Z0 => UQVN_N184, A0 => A0, A1 => B1);
UQVB_B222 : AND2
	PORT MAP (Z0 => UQVN_N183, A0 => UQVN_N206, A1 => B1);
UQVB_B223 : OR3
	PORT MAP (Z0 => UQVN_N186, A0 => UQVN_N184, A1 => UQVN_N183, A2 => UQVN_N185);
UQVB_B224 : INV
	PORT MAP (ZN0 => UQVN_N208, A0 => B2);
UQVB_B225 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B226 : INV
	PORT MAP (ZN0 => UQVN_N205, A0 => A2);
UQVB_B227 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N198);
UQVB_B228 : AND4
	PORT MAP (Z0 => UQVN_N197, A0 => UQVN_N203, A1 => B0, A2 => B1, 
	A3 => UQVN_N208);
UQVB_B229 : AND3
	PORT MAP (Z0 => UQVN_N196, A0 => A1, A1 => UQVN_N207, A2 => B2);
UQVB_B230 : AND4
	PORT MAP (Z0 => UQVN_N195, A0 => UQVN_N203, A1 => UQVN_N204, A2 => B0, 
	A3 => UQVN_N208);
UQVB_B231 : AND3
	PORT MAP (Z0 => UQVN_N194, A0 => UQVN_N206, A1 => UQVN_N207, A2 => B2);
UQVB_B232 : AND3
	PORT MAP (Z0 => UQVN_N202, A0 => A0, A1 => A1, A2 => B2);
UQVB_B233 : AND3
	PORT MAP (Z0 => UQVN_N201, A0 => A1, A1 => UQVN_N206, A2 => B2);
UQVB_B234 : AND3
	PORT MAP (Z0 => UQVN_N200, A0 => UQVN_N204, A1 => B1, A2 => UQVN_N208);
UQVB_B235 : AND3
	PORT MAP (Z0 => UQVN_N199, A0 => A0, A1 => UQVN_N207, A2 => B2);
UQVB_B236 : OR8
	PORT MAP (Z0 => UQVN_N198, A0 => UQVN_N202, A1 => UQVN_N201, A2 => UQVN_N200, 
	A3 => UQVN_N199, A4 => UQVN_N197, A5 => UQVN_N196, A6 => UQVN_N195, 
	A7 => UQVN_N194);
UQVB_B237 : XOR2
	PORT MAP (Z0 => Z15, A0 => A15, A1 => UQVN_N212);
UQVB_B238 : AND2
	PORT MAP (Z0 => UQVN_N211, A0 => UQVN_N217, A1 => UQVN_N221);
UQVB_B239 : AND2
	PORT MAP (Z0 => UQVN_N210, A0 => B15, A1 => UQVN_N209);
UQVB_B240 : OR2
	PORT MAP (Z0 => UQVN_N212, A0 => UQVN_N210, A1 => UQVN_N211);
UQVB_B241 : INV
	PORT MAP (ZN0 => UQVN_N213, A0 => A15);
UQVB_B242 : INV
	PORT MAP (ZN0 => UQVN_N217, A0 => B15);
UQVB_B243 : INV
	PORT MAP (ZN0 => UQVN_N209, A0 => UQVN_N221);
UQVB_B244 : AND2
	PORT MAP (Z0 => UQVN_N214, A0 => UQVN_N221, A1 => B15);
UQVB_B245 : AND2
	PORT MAP (Z0 => UQVN_N215, A0 => UQVN_N221, A1 => UQVN_N213);
UQVB_B246 : AND2
	PORT MAP (Z0 => UQVN_N216, A0 => B15, A1 => UQVN_N213);
UQVB_B247 : OR3
	PORT MAP (Z0 => BO, A0 => UQVN_N214, A1 => UQVN_N215, A2 => UQVN_N216);
END lattice_arch;
-- VHDL netlist for SUBH2
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH2 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBH2;


ARCHITECTURE lattice_arch OF SUBH2 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N12, A1 => B0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N14);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N13, A1 => UQVN_N12, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N12, A1 => B1, A2 => B0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N13, A1 => B1);
UQVB_B6 : OR3
	PORT MAP (Z0 => BO, A0 => UQVN_N3, A1 => UQVN_N5, A2 => UQVN_N4);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => B0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => B1);
UQVB_B10 : OR6
	PORT MAP (Z0 => Z1, A0 => UQVN_N6, A1 => UQVN_N8, A2 => UQVN_N7, 
	A3 => UQVN_N9, A4 => UQVN_N10, A5 => UQVN_N11);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N13, A1 => B1, A2 => A0);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N13, A1 => B1, A2 => UQVN_N14);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N15, A2 => A0);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => A1, A1 => UQVN_N15, A2 => UQVN_N14);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N13, A1 => UQVN_N15, A2 => UQVN_N12, 
	A3 => B0);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A1, A1 => B1, A2 => UQVN_N12, 
	A3 => B0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => A0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => A1);
END lattice_arch;
-- VHDL netlist for SUBH3
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH3 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBH3;


ARCHITECTURE lattice_arch OF SUBH3 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26 : std_logic;


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


BEGIN

UQVB_B1 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => B1);
UQVB_B2 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => A0);
UQVB_B3 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N4);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N21, A1 => B0, A2 => UQVN_N25);
UQVB_B5 : AND4
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N21, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B6 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => UQVN_N22, A1 => B1, A2 => B2);
UQVB_B7 : AND4
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N21, A1 => UQVN_N23, A2 => B0, 
	A3 => B1);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N23, A1 => B2);
UQVB_B9 : AND4
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N21, A1 => UQVN_N22, A2 => UQVN_N23, 
	A3 => B0);
UQVB_B10 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N22, A1 => UQVN_N23, A2 => B1);
UQVB_B11 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N21, A1 => UQVN_N22, A2 => B0, 
	A3 => B2);
UQVB_B12 : OR7
	PORT MAP (Z0 => BO, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N6, 
	A3 => UQVN_N5, A4 => UQVN_N9, A5 => UQVN_N10, A6 => UQVN_N11);
UQVB_B13 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => B0);
UQVB_B14 : INV
	PORT MAP (ZN0 => UQVN_N22, A0 => A1);
UQVB_B15 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => A0, A1 => B1);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N24, A1 => B1);
UQVB_B17 : OR3
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N2, A1 => UQVN_N1, A2 => UQVN_N3);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => B2);
UQVB_B19 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => A2);
UQVB_B21 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N16);
UQVB_B22 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N21, A1 => B0, A2 => B1, 
	A3 => UQVN_N26);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => A1, A1 => UQVN_N25, A2 => B2);
UQVB_B24 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N21, A1 => UQVN_N22, A2 => B0, 
	A3 => UQVN_N26);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N24, A1 => UQVN_N25, A2 => B2);
UQVB_B26 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => A0, A1 => A1, A2 => B2);
UQVB_B27 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => A1, A1 => UQVN_N24, A2 => B2);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N22, A1 => B1, A2 => UQVN_N26);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => A0, A1 => UQVN_N25, A2 => B2);
UQVB_B30 : OR8
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N20, A1 => UQVN_N19, A2 => UQVN_N18, 
	A3 => UQVN_N17, A4 => UQVN_N15, A5 => UQVN_N14, A6 => UQVN_N13, 
	A7 => UQVN_N12);
END lattice_arch;
-- VHDL netlist for SUBH4
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH4 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBH4;


ARCHITECTURE lattice_arch OF SUBH4 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N12, A1 => B0);
UQVB_B2 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => A0, A1 => UQVN_N14);
UQVB_B3 : AND3
	PORT MAP (Z0 => UQVN_N3, A0 => UQVN_N13, A1 => UQVN_N12, A2 => B0);
UQVB_B4 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N12, A1 => B1, A2 => B0);
UQVB_B5 : AND2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N13, A1 => B1);
UQVB_B6 : OR3
	PORT MAP (Z0 => UQVN_N38, A0 => UQVN_N3, A1 => UQVN_N5, A2 => UQVN_N4);
UQVB_B7 : OR2
	PORT MAP (Z0 => Z0, A0 => UQVN_N2, A1 => UQVN_N1);
UQVB_B8 : INV
	PORT MAP (ZN0 => UQVN_N14, A0 => B0);
UQVB_B9 : INV
	PORT MAP (ZN0 => UQVN_N15, A0 => B1);
UQVB_B10 : OR6
	PORT MAP (Z0 => Z1, A0 => UQVN_N6, A1 => UQVN_N8, A2 => UQVN_N7, 
	A3 => UQVN_N9, A4 => UQVN_N10, A5 => UQVN_N11);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N13, A1 => B1, A2 => A0);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => UQVN_N13, A1 => B1, A2 => UQVN_N14);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => A1, A1 => UQVN_N15, A2 => A0);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => A1, A1 => UQVN_N15, A2 => UQVN_N14);
UQVB_B15 : AND4
	PORT MAP (Z0 => UQVN_N10, A0 => UQVN_N13, A1 => UQVN_N15, A2 => UQVN_N12, 
	A3 => B0);
UQVB_B16 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => A1, A1 => B1, A2 => UQVN_N12, 
	A3 => B0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N12, A0 => A0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N13, A0 => A1);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N37, A0 => UQVN_N38);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N38, A1 => UQVN_N34, A2 => UQVN_N33);
UQVB_B21 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N38, A1 => UQVN_N34, A2 => B2);
UQVB_B22 : AND3
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N38, A1 => UQVN_N33, A2 => B3);
UQVB_B23 : AND3
	PORT MAP (Z0 => UQVN_N19, A0 => UQVN_N38, A1 => B3, A2 => B2);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N34, A1 => UQVN_N33, A2 => B2);
UQVB_B25 : AND3
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N33, A1 => B3, A2 => B2);
UQVB_B26 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => UQVN_N34, A1 => B3);
UQVB_B27 : OR7
	PORT MAP (Z0 => BO, A0 => UQVN_N18, A1 => UQVN_N17, A2 => UQVN_N16, 
	A3 => UQVN_N19, A4 => UQVN_N20, A5 => UQVN_N22, A6 => UQVN_N21);
UQVB_B28 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => A2, A1 => B3, A2 => UQVN_N37);
UQVB_B29 : AND3
	PORT MAP (Z0 => UQVN_N24, A0 => B3, A1 => UQVN_N35, A2 => UQVN_N37);
UQVB_B30 : AND3
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N33, A1 => UQVN_N36, A2 => UQVN_N38);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N36, A1 => B2, A2 => UQVN_N38);
UQVB_B32 : AND3
	PORT MAP (Z0 => UQVN_N27, A0 => A2, A1 => B3, A2 => UQVN_N35);
UQVB_B33 : AND3
	PORT MAP (Z0 => UQVN_N28, A0 => UQVN_N33, A1 => UQVN_N36, A2 => B2);
UQVB_B34 : OR6
	PORT MAP (Z0 => UQVN_N29, A0 => UQVN_N23, A1 => UQVN_N24, A2 => UQVN_N25, 
	A3 => UQVN_N26, A4 => UQVN_N27, A5 => UQVN_N28);
UQVB_B35 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N29);
UQVB_B36 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => B2);
UQVB_B37 : INV
	PORT MAP (ZN0 => UQVN_N36, A0 => B3);
UQVB_B38 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => A3);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => A2);
UQVB_B40 : XOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N30);
UQVB_B41 : OR2
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N31, A1 => UQVN_N32);
UQVB_B42 : AND2
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N35, A1 => UQVN_N38);
UQVB_B43 : AND2
	PORT MAP (Z0 => UQVN_N32, A0 => UQVN_N37, A1 => B2);
END lattice_arch;
-- VHDL netlist for SUBH8
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH8 IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBH8;


ARCHITECTURE lattice_arch OF SUBH8 IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 G1, G2, G3, G4,
	 G5, G6, G7, P1,
	 P2, P3, P4, P5,
	 P6, P7 : std_logic;


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND9
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND9 use  entity  lat_vhd.AND9(lattice_arch);


  COMPONENT OR5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR5 use  entity  lat_vhd.OR5(lattice_arch);


  COMPONENT AND7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND7 use  entity  lat_vhd.AND7(lattice_arch);


  COMPONENT OR4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR4 use  entity  lat_vhd.OR4(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT AND6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND6 use  entity  lat_vhd.AND6(lattice_arch);


  COMPONENT AND5
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND5 use  entity  lat_vhd.AND5(lattice_arch);


  COMPONENT AND8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND8 use  entity  lat_vhd.AND8(lattice_arch);


BEGIN

UQVB_B1 : XOR2
	PORT MAP (Z0 => P7, A0 => A7, A1 => B7);
UQVB_B2 : XOR2
	PORT MAP (Z0 => P6, A0 => A6, A1 => B6);
UQVB_B3 : XOR2
	PORT MAP (Z0 => P5, A0 => A5, A1 => B5);
UQVB_B4 : XOR2
	PORT MAP (Z0 => P4, A0 => A4, A1 => B4);
UQVB_B5 : XOR2
	PORT MAP (Z0 => P3, A0 => A3, A1 => B3);
UQVB_B6 : XOR2
	PORT MAP (Z0 => P2, A0 => A2, A1 => B2);
UQVB_B7 : XOR2
	PORT MAP (Z0 => P1, A0 => A1, A1 => B1);
UQVB_B8 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B9 : AND2
	PORT MAP (Z0 => G7, A0 => UQVN_N9, A1 => B7);
UQVB_B10 : AND2
	PORT MAP (Z0 => G6, A0 => UQVN_N8, A1 => B6);
UQVB_B11 : AND2
	PORT MAP (Z0 => G5, A0 => UQVN_N7, A1 => B5);
UQVB_B12 : AND2
	PORT MAP (Z0 => G4, A0 => UQVN_N6, A1 => B4);
UQVB_B13 : AND2
	PORT MAP (Z0 => G3, A0 => UQVN_N5, A1 => B3);
UQVB_B14 : AND2
	PORT MAP (Z0 => G2, A0 => UQVN_N4, A1 => B2);
UQVB_B15 : AND2
	PORT MAP (Z0 => G1, A0 => UQVN_N3, A1 => B1);
UQVB_B16 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => UQVN_N2, A1 => B0);
UQVB_B17 : INV
	PORT MAP (ZN0 => UQVN_N2, A0 => A0);
UQVB_B18 : INV
	PORT MAP (ZN0 => UQVN_N3, A0 => A1);
UQVB_B19 : INV
	PORT MAP (ZN0 => UQVN_N4, A0 => A2);
UQVB_B20 : INV
	PORT MAP (ZN0 => UQVN_N5, A0 => A3);
UQVB_B21 : INV
	PORT MAP (ZN0 => UQVN_N6, A0 => A4);
UQVB_B22 : INV
	PORT MAP (ZN0 => UQVN_N7, A0 => A5);
UQVB_B23 : INV
	PORT MAP (ZN0 => UQVN_N8, A0 => A6);
UQVB_B24 : INV
	PORT MAP (ZN0 => UQVN_N9, A0 => A7);
UQVB_B25 : LXOR2
	PORT MAP (Z0 => Z1, A0 => P1, A1 => UQVN_N1);
UQVB_B26 : AND9
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N24, A1 => B0, A2 => UQVN_N23, 
	A3 => UQVN_N35, A4 => UQVN_N34, A5 => UQVN_N33, A6 => UQVN_N32, 
	A7 => UQVN_N30, A8 => UQVN_N17);
UQVB_B27 : OR5
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N12, A1 => UQVN_N11, A2 => UQVN_N13, 
	A3 => UQVN_N14, A4 => G4);
UQVB_B28 : LXOR2
	PORT MAP (Z0 => Z5, A0 => UQVN_N15, A1 => P5);
UQVB_B29 : AND7
	PORT MAP (Z0 => UQVN_N36, A0 => G1, A1 => UQVN_N35, A2 => UQVN_N34, 
	A3 => UQVN_N33, A4 => UQVN_N32, A5 => UQVN_N30, A6 => UQVN_N17);
UQVB_B30 : OR4
	PORT MAP (Z0 => UQVN_N43, A0 => UQVN_N39, A1 => UQVN_N42, A2 => UQVN_N41, 
	A3 => G7);
UQVB_B31 : AND3
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N25, A1 => B0, A2 => UQVN_N26);
UQVB_B32 : OR2
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N18, A1 => G1);
UQVB_B33 : LXOR2
	PORT MAP (Z0 => Z2, A0 => UQVN_N16, A1 => P2);
UQVB_B34 : OR4
	PORT MAP (Z0 => UQVN_N44, A0 => UQVN_N37, A1 => UQVN_N36, A2 => UQVN_N38, 
	A3 => UQVN_N40);
UQVB_B35 : OR3
	PORT MAP (Z0 => UQVN_N20, A0 => UQVN_N22, A1 => UQVN_N19, A2 => G2);
UQVB_B36 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => G1, A1 => UQVN_N21);
UQVB_B37 : LXOR2
	PORT MAP (Z0 => Z3, A0 => UQVN_N20, A1 => P3);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => UQVN_N29, A1 => B0, A2 => UQVN_N31, 
	A3 => UQVN_N21);
UQVB_B39 : INV
	PORT MAP (ZN0 => UQVN_N17, A0 => P7);
UQVB_B40 : INV
	PORT MAP (ZN0 => UQVN_N30, A0 => P6);
UQVB_B41 : INV
	PORT MAP (ZN0 => UQVN_N32, A0 => P5);
UQVB_B42 : INV
	PORT MAP (ZN0 => UQVN_N33, A0 => P4);
UQVB_B43 : INV
	PORT MAP (ZN0 => UQVN_N34, A0 => P3);
UQVB_B44 : INV
	PORT MAP (ZN0 => UQVN_N35, A0 => P2);
UQVB_B45 : AND6
	PORT MAP (Z0 => UQVN_N38, A0 => G2, A1 => UQVN_N34, A2 => UQVN_N33, 
	A3 => UQVN_N32, A4 => UQVN_N30, A5 => UQVN_N17);
UQVB_B46 : INV
	PORT MAP (ZN0 => UQVN_N23, A0 => P1);
UQVB_B47 : INV
	PORT MAP (ZN0 => UQVN_N24, A0 => A0);
UQVB_B48 : INV
	PORT MAP (ZN0 => UQVN_N25, A0 => A0);
UQVB_B49 : INV
	PORT MAP (ZN0 => UQVN_N26, A0 => P1);
UQVB_B50 : INV
	PORT MAP (ZN0 => UQVN_N45, A0 => P4);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N46, A0 => P3);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N10, A0 => P2);
UQVB_B53 : INV
	PORT MAP (ZN0 => UQVN_N28, A0 => P1);
UQVB_B54 : INV
	PORT MAP (ZN0 => UQVN_N27, A0 => A0);
UQVB_B55 : INV
	PORT MAP (ZN0 => UQVN_N21, A0 => P2);
UQVB_B56 : INV
	PORT MAP (ZN0 => UQVN_N31, A0 => P1);
UQVB_B57 : INV
	PORT MAP (ZN0 => UQVN_N29, A0 => A0);
UQVB_B58 : AND5
	PORT MAP (Z0 => UQVN_N40, A0 => G3, A1 => UQVN_N33, A2 => UQVN_N32, 
	A3 => UQVN_N30, A4 => UQVN_N17);
UQVB_B59 : AND2
	PORT MAP (Z0 => UQVN_N41, A0 => G6, A1 => UQVN_N17);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N42, A0 => G5, A1 => UQVN_N30, A2 => UQVN_N17);
UQVB_B61 : AND4
	PORT MAP (Z0 => UQVN_N39, A0 => G4, A1 => UQVN_N32, A2 => UQVN_N30, 
	A3 => UQVN_N17);
UQVB_B62 : OR2
	PORT MAP (Z0 => BO, A0 => UQVN_N44, A1 => UQVN_N43);
UQVB_B63 : AND6
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N27, A1 => B0, A2 => UQVN_N28, 
	A3 => UQVN_N10, A4 => UQVN_N46, A5 => UQVN_N45);
UQVB_B64 : AND4
	PORT MAP (Z0 => UQVN_N11, A0 => G1, A1 => UQVN_N10, A2 => UQVN_N46, 
	A3 => UQVN_N45);
UQVB_B65 : AND3
	PORT MAP (Z0 => UQVN_N13, A0 => G2, A1 => UQVN_N46, A2 => UQVN_N45);
UQVB_B66 : AND2
	PORT MAP (Z0 => UQVN_N14, A0 => G3, A1 => UQVN_N45);
UQVB_B67 : AND3
	PORT MAP (Z0 => UQVN_N50, A0 => G3, A1 => UQVN_N56, A2 => UQVN_N57);
UQVB_B68 : AND4
	PORT MAP (Z0 => UQVN_N51, A0 => G2, A1 => UQVN_N55, A2 => UQVN_N56, 
	A3 => UQVN_N57);
UQVB_B69 : AND5
	PORT MAP (Z0 => UQVN_N48, A0 => G1, A1 => UQVN_N54, A2 => UQVN_N55, 
	A3 => UQVN_N56, A4 => UQVN_N57);
UQVB_B70 : AND2
	PORT MAP (Z0 => UQVN_N49, A0 => G4, A1 => UQVN_N57);
UQVB_B71 : OR3
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N50, A1 => UQVN_N49, A2 => G5);
UQVB_B72 : OR3
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N58, A1 => UQVN_N48, A2 => UQVN_N51);
UQVB_B73 : OR2
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N53, A1 => UQVN_N52);
UQVB_B74 : LXOR2
	PORT MAP (Z0 => Z6, A0 => UQVN_N47, A1 => P6);
UQVB_B75 : AND7
	PORT MAP (Z0 => UQVN_N58, A0 => UQVN_N70, A1 => B0, A2 => UQVN_N69, 
	A3 => UQVN_N54, A4 => UQVN_N55, A5 => UQVN_N56, A6 => UQVN_N57);
UQVB_B76 : AND5
	PORT MAP (Z0 => UQVN_N64, A0 => UQVN_N71, A1 => B0, A2 => UQVN_N72, 
	A3 => UQVN_N63, A4 => UQVN_N62);
UQVB_B77 : AND3
	PORT MAP (Z0 => UQVN_N59, A0 => G1, A1 => UQVN_N63, A2 => UQVN_N62);
UQVB_B78 : AND2
	PORT MAP (Z0 => UQVN_N60, A0 => G2, A1 => UQVN_N62);
UQVB_B79 : OR4
	PORT MAP (Z0 => UQVN_N61, A0 => UQVN_N64, A1 => UQVN_N59, A2 => UQVN_N60, 
	A3 => G3);
UQVB_B80 : LXOR2
	PORT MAP (Z0 => Z4, A0 => UQVN_N61, A1 => P4);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N75, A0 => P6);
UQVB_B82 : INV
	PORT MAP (ZN0 => UQVN_N74, A0 => P5);
UQVB_B83 : INV
	PORT MAP (ZN0 => UQVN_N73, A0 => P4);
UQVB_B84 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => P3);
UQVB_B85 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => P1);
UQVB_B86 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => A0);
UQVB_B87 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => P2);
UQVB_B88 : INV
	PORT MAP (ZN0 => UQVN_N54, A0 => P2);
UQVB_B89 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => P1);
UQVB_B90 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => A0);
UQVB_B91 : INV
	PORT MAP (ZN0 => UQVN_N55, A0 => P3);
UQVB_B92 : INV
	PORT MAP (ZN0 => UQVN_N56, A0 => P4);
UQVB_B93 : INV
	PORT MAP (ZN0 => UQVN_N57, A0 => P5);
UQVB_B94 : INV
	PORT MAP (ZN0 => UQVN_N63, A0 => P2);
UQVB_B95 : INV
	PORT MAP (ZN0 => UQVN_N62, A0 => P3);
UQVB_B96 : INV
	PORT MAP (ZN0 => UQVN_N72, A0 => P1);
UQVB_B97 : INV
	PORT MAP (ZN0 => UQVN_N71, A0 => A0);
UQVB_B98 : OR2
	PORT MAP (Z0 => UQVN_N84, A0 => UQVN_N77, A1 => UQVN_N76);
UQVB_B99 : AND2
	PORT MAP (Z0 => UQVN_N83, A0 => G5, A1 => UQVN_N75);
UQVB_B100 : AND3
	PORT MAP (Z0 => UQVN_N81, A0 => G4, A1 => UQVN_N74, A2 => UQVN_N75);
UQVB_B101 : AND4
	PORT MAP (Z0 => UQVN_N82, A0 => G3, A1 => UQVN_N73, A2 => UQVN_N74, 
	A3 => UQVN_N75);
UQVB_B102 : AND5
	PORT MAP (Z0 => UQVN_N80, A0 => G2, A1 => UQVN_N68, A2 => UQVN_N73, 
	A3 => UQVN_N74, A4 => UQVN_N75);
UQVB_B103 : AND6
	PORT MAP (Z0 => UQVN_N78, A0 => G1, A1 => UQVN_N67, A2 => UQVN_N68, 
	A3 => UQVN_N73, A4 => UQVN_N74, A5 => UQVN_N75);
UQVB_B104 : AND8
	PORT MAP (Z0 => UQVN_N79, A0 => UQVN_N66, A1 => B0, A2 => UQVN_N65, 
	A3 => UQVN_N67, A4 => UQVN_N68, A5 => UQVN_N73, A6 => UQVN_N74, 
	A7 => UQVN_N75);
UQVB_B105 : OR4
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N79, A1 => UQVN_N78, A2 => UQVN_N80, 
	A3 => UQVN_N82);
UQVB_B106 : OR3
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N81, A1 => UQVN_N83, A2 => G6);
UQVB_B107 : LXOR2
	PORT MAP (Z0 => Z7, A0 => UQVN_N84, A1 => P7);
END lattice_arch;
-- VHDL netlist for SUBH8A
-- Date: 15.5.95 13.47.13

LIBRARY IEEE;
LIBRARY lat_vhd;
USE lat_vhd.vhd_pkg.all;
USE IEEE.std_logic_1164.all;
USE work.all;

ENTITY SUBH8A IS 
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        B0 : IN std_logic;
        B1 : IN std_logic;
        B2 : IN std_logic;
        B3 : IN std_logic;
        B4 : IN std_logic;
        B5 : IN std_logic;
        B6 : IN std_logic;
        B7 : IN std_logic;
        Z0 : OUT std_logic;
        Z1 : OUT std_logic;
        Z2 : OUT std_logic;
        Z3 : OUT std_logic;
        Z4 : OUT std_logic;
        Z5 : OUT std_logic;
        Z6 : OUT std_logic;
        Z7 : OUT std_logic;
        BO : OUT std_logic
    );
END SUBH8A;


ARCHITECTURE lattice_arch OF SUBH8A IS
SIGNAL  UQVN_N1, UQVN_N2, UQVN_N3, UQVN_N4,
	 UQVN_N5, UQVN_N6, UQVN_N7, UQVN_N8,
	 UQVN_N9, UQVN_N10, UQVN_N11, UQVN_N12,
	 UQVN_N13, UQVN_N14, UQVN_N15, UQVN_N16,
	 UQVN_N17, UQVN_N18, UQVN_N19, UQVN_N20,
	 UQVN_N21, UQVN_N22, UQVN_N23, UQVN_N24,
	 UQVN_N25, UQVN_N26, UQVN_N27, UQVN_N28,
	 UQVN_N29, UQVN_N30, UQVN_N31, UQVN_N32,
	 UQVN_N33, UQVN_N34, UQVN_N35, UQVN_N36,
	 UQVN_N37, UQVN_N38, UQVN_N39, UQVN_N40,
	 UQVN_N41, UQVN_N42, UQVN_N43, UQVN_N44,
	 UQVN_N45, UQVN_N46, UQVN_N47, UQVN_N48,
	 UQVN_N49, UQVN_N50, UQVN_N51, UQVN_N52,
	 UQVN_N53, UQVN_N54, UQVN_N55, UQVN_N56,
	 UQVN_N57, UQVN_N58, UQVN_N59, UQVN_N60,
	 UQVN_N61, UQVN_N62, UQVN_N63, UQVN_N64,
	 UQVN_N65, UQVN_N66, UQVN_N67, UQVN_N68,
	 UQVN_N69, UQVN_N70, UQVN_N71, UQVN_N72,
	 UQVN_N73, UQVN_N74, UQVN_N75, UQVN_N76,
	 UQVN_N77, UQVN_N78, UQVN_N79, UQVN_N80,
	 UQVN_N81, UQVN_N82, UQVN_N83, UQVN_N84,
	 UQVN_N85, UQVN_N86, UQVN_N87, UQVN_N88,
	 UQVN_N89, UQVN_N90, UQVN_N91, UQVN_N92,
	 UQVN_N93, G012, G345, P345 : std_logic;


  COMPONENT AND2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND2 use  entity  lat_vhd.AND2(lattice_arch);


  COMPONENT OR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR2 use  entity  lat_vhd.OR2(lattice_arch);


  COMPONENT INV
    PORT (
        A0 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: INV use  entity  lat_vhd.INV(lattice_arch);


  COMPONENT LXOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: LXOR2 use  entity  lat_vhd.LXOR2(lattice_arch);


  COMPONENT AND3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND3 use  entity  lat_vhd.AND3(lattice_arch);


  COMPONENT OR6
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR6 use  entity  lat_vhd.OR6(lattice_arch);


  COMPONENT AND4
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: AND4 use  entity  lat_vhd.AND4(lattice_arch);


  COMPONENT OR7
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR7 use  entity  lat_vhd.OR7(lattice_arch);


  COMPONENT NOR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        ZN0 : OUT std_logic
    );
  END COMPONENT;

for all: NOR3 use  entity  lat_vhd.NOR3(lattice_arch);


  COMPONENT OR12
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        A8 : IN std_logic;
        A9 : IN std_logic;
        A10 : IN std_logic;
        A11 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR12 use  entity  lat_vhd.OR12(lattice_arch);


  COMPONENT OR3
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR3 use  entity  lat_vhd.OR3(lattice_arch);


  COMPONENT XOR2
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: XOR2 use  entity  lat_vhd.XOR2(lattice_arch);


  COMPONENT OR8
    PORT (
        A0 : IN std_logic;
        A1 : IN std_logic;
        A2 : IN std_logic;
        A3 : IN std_logic;
        A4 : IN std_logic;
        A5 : IN std_logic;
        A6 : IN std_logic;
        A7 : IN std_logic;
        Z0 : OUT std_logic
    );
  END COMPONENT;

for all: OR8 use  entity  lat_vhd.OR8(lattice_arch);


BEGIN

UQVB_B1 : AND2
	PORT MAP (Z0 => UQVN_N1, A0 => P345, A1 => G012);
UQVB_B2 : OR2
	PORT MAP (Z0 => UQVN_N93, A0 => G345, A1 => UQVN_N1);
UQVB_B3 : INV
	PORT MAP (ZN0 => UQVN_N44, A0 => G012);
UQVB_B4 : INV
	PORT MAP (ZN0 => UQVN_N42, A0 => B4);
UQVB_B5 : INV
	PORT MAP (ZN0 => UQVN_N43, A0 => B5);
UQVB_B6 : INV
	PORT MAP (ZN0 => UQVN_N38, A0 => A3);
UQVB_B7 : AND2
	PORT MAP (Z0 => UQVN_N2, A0 => UQVN_N41, A1 => G012);
UQVB_B8 : AND2
	PORT MAP (Z0 => UQVN_N3, A0 => B3, A1 => UQVN_N44);
UQVB_B9 : OR2
	PORT MAP (Z0 => UQVN_N4, A0 => UQVN_N2, A1 => UQVN_N3);
UQVB_B10 : LXOR2
	PORT MAP (Z0 => Z3, A0 => A3, A1 => UQVN_N4);
UQVB_B11 : AND3
	PORT MAP (Z0 => UQVN_N10, A0 => A3, A1 => B4, A2 => UQVN_N41);
UQVB_B12 : AND3
	PORT MAP (Z0 => UQVN_N6, A0 => UQVN_N42, A1 => B3, A2 => G012);
UQVB_B13 : AND3
	PORT MAP (Z0 => UQVN_N5, A0 => UQVN_N38, A1 => UQVN_N42, A2 => G012);
UQVB_B14 : AND3
	PORT MAP (Z0 => UQVN_N7, A0 => B4, A1 => UQVN_N41, A2 => UQVN_N44);
UQVB_B15 : AND3
	PORT MAP (Z0 => UQVN_N8, A0 => A3, A1 => B4, A2 => UQVN_N44);
UQVB_B16 : OR6
	PORT MAP (Z0 => UQVN_N11, A0 => UQVN_N8, A1 => UQVN_N7, A2 => UQVN_N5, 
	A3 => UQVN_N6, A4 => UQVN_N10, A5 => UQVN_N9);
UQVB_B17 : LXOR2
	PORT MAP (Z0 => Z4, A0 => A4, A1 => UQVN_N11);
UQVB_B18 : AND3
	PORT MAP (Z0 => UQVN_N9, A0 => UQVN_N38, A1 => UQVN_N42, A2 => B3);
UQVB_B19 : AND4
	PORT MAP (Z0 => UQVN_N15, A0 => UQVN_N38, A1 => B3, A2 => B4, 
	A3 => B5);
UQVB_B20 : AND3
	PORT MAP (Z0 => UQVN_N14, A0 => UQVN_N39, A1 => B4, A2 => B5);
UQVB_B21 : AND4
	PORT MAP (Z0 => UQVN_N13, A0 => UQVN_N38, A1 => UQVN_N40, A2 => B3, 
	A3 => B4);
UQVB_B22 : AND2
	PORT MAP (Z0 => UQVN_N12, A0 => UQVN_N40, A1 => B5);
UQVB_B23 : AND4
	PORT MAP (Z0 => UQVN_N16, A0 => UQVN_N38, A1 => UQVN_N39, A2 => B3, 
	A3 => B5);
UQVB_B24 : AND3
	PORT MAP (Z0 => UQVN_N17, A0 => UQVN_N39, A1 => UQVN_N40, A2 => B4);
UQVB_B25 : AND4
	PORT MAP (Z0 => UQVN_N18, A0 => UQVN_N38, A1 => UQVN_N39, A2 => UQVN_N40, 
	A3 => B3);
UQVB_B26 : OR7
	PORT MAP (Z0 => G345, A0 => UQVN_N15, A1 => UQVN_N14, A2 => UQVN_N13, 
	A3 => UQVN_N12, A4 => UQVN_N16, A5 => UQVN_N17, A6 => UQVN_N18);
UQVB_B27 : AND2
	PORT MAP (Z0 => UQVN_N21, A0 => A3, A1 => UQVN_N41);
UQVB_B28 : AND2
	PORT MAP (Z0 => UQVN_N19, A0 => A4, A1 => UQVN_N42);
UQVB_B29 : AND2
	PORT MAP (Z0 => UQVN_N20, A0 => A5, A1 => UQVN_N43);
UQVB_B30 : NOR3
	PORT MAP (ZN0 => P345, A0 => UQVN_N21, A1 => UQVN_N19, A2 => UQVN_N20);
UQVB_B31 : INV
	PORT MAP (ZN0 => UQVN_N41, A0 => B3);
UQVB_B32 : INV
	PORT MAP (ZN0 => UQVN_N39, A0 => A4);
UQVB_B33 : INV
	PORT MAP (ZN0 => UQVN_N40, A0 => A5);
UQVB_B34 : LXOR2
	PORT MAP (Z0 => Z5, A0 => A5, A1 => UQVN_N35);
UQVB_B35 : AND4
	PORT MAP (Z0 => UQVN_N34, A0 => A3, A1 => A4, A2 => B5, 
	A3 => UQVN_N44);
UQVB_B36 : AND4
	PORT MAP (Z0 => UQVN_N36, A0 => UQVN_N38, A1 => UQVN_N39, A2 => UQVN_N43, 
	A3 => G012);
UQVB_B37 : AND4
	PORT MAP (Z0 => UQVN_N33, A0 => A3, A1 => A4, A2 => UQVN_N41, 
	A3 => B5);
UQVB_B38 : AND4
	PORT MAP (Z0 => UQVN_N32, A0 => A4, A1 => UQVN_N41, A2 => B5, 
	A3 => UQVN_N44);
UQVB_B39 : AND4
	PORT MAP (Z0 => UQVN_N31, A0 => UQVN_N38, A1 => UQVN_N39, A2 => B3, 
	A3 => UQVN_N43);
UQVB_B40 : AND4
	PORT MAP (Z0 => UQVN_N30, A0 => UQVN_N39, A1 => B3, A2 => UQVN_N43, 
	A3 => G012);
UQVB_B41 : AND4
	PORT MAP (Z0 => UQVN_N29, A0 => A3, A1 => UQVN_N42, A2 => B5, 
	A3 => UQVN_N44);
UQVB_B42 : AND4
	PORT MAP (Z0 => UQVN_N28, A0 => A3, A1 => UQVN_N41, A2 => UQVN_N42, 
	A3 => B5);
UQVB_B43 : AND4
	PORT MAP (Z0 => UQVN_N27, A0 => UQVN_N41, A1 => UQVN_N42, A2 => B5, 
	A3 => UQVN_N44);
UQVB_B44 : AND3
	PORT MAP (Z0 => UQVN_N26, A0 => UQVN_N39, A1 => UQVN_N43, A2 => B4);
UQVB_B45 : AND4
	PORT MAP (Z0 => UQVN_N25, A0 => UQVN_N38, A1 => B4, A2 => UQVN_N43, 
	A3 => G012);
UQVB_B46 : AND4
	PORT MAP (Z0 => UQVN_N24, A0 => UQVN_N38, A1 => B3, A2 => B4, 
	A3 => UQVN_N43);
UQVB_B47 : AND3
	PORT MAP (Z0 => UQVN_N23, A0 => A4, A1 => UQVN_N42, A2 => B5);
UQVB_B48 : AND4
	PORT MAP (Z0 => UQVN_N22, A0 => B3, A1 => B4, A2 => UQVN_N43, 
	A3 => G012);
UQVB_B49 : OR12
	PORT MAP (Z0 => UQVN_N37, A0 => UQVN_N33, A1 => UQVN_N32, A2 => UQVN_N31, 
	A3 => UQVN_N30, A4 => UQVN_N29, A5 => UQVN_N28, A6 => UQVN_N27, 
	A7 => UQVN_N26, A8 => UQVN_N25, A9 => UQVN_N24, A10 => UQVN_N23, 
	A11 => UQVN_N22);
UQVB_B50 : OR3
	PORT MAP (Z0 => UQVN_N35, A0 => UQVN_N34, A1 => UQVN_N36, A2 => UQVN_N37);
UQVB_B51 : INV
	PORT MAP (ZN0 => UQVN_N69, A0 => B1);
UQVB_B52 : INV
	PORT MAP (ZN0 => UQVN_N65, A0 => A0);
UQVB_B53 : LXOR2
	PORT MAP (Z0 => Z1, A0 => A1, A1 => UQVN_N48);
UQVB_B54 : AND3
	PORT MAP (Z0 => UQVN_N47, A0 => UQVN_N65, A1 => B0, A2 => UQVN_N69);
UQVB_B55 : AND4
	PORT MAP (Z0 => UQVN_N52, A0 => UQVN_N65, A1 => B0, A2 => B1, 
	A3 => B2);
UQVB_B56 : AND3
	PORT MAP (Z0 => UQVN_N51, A0 => UQVN_N66, A1 => B1, A2 => B2);
UQVB_B57 : AND4
	PORT MAP (Z0 => UQVN_N50, A0 => UQVN_N65, A1 => UQVN_N67, A2 => B0, 
	A3 => B1);
UQVB_B58 : AND2
	PORT MAP (Z0 => UQVN_N49, A0 => UQVN_N67, A1 => B2);
UQVB_B59 : AND4
	PORT MAP (Z0 => UQVN_N53, A0 => UQVN_N65, A1 => UQVN_N66, A2 => UQVN_N67, 
	A3 => B0);
UQVB_B60 : AND3
	PORT MAP (Z0 => UQVN_N54, A0 => UQVN_N66, A1 => UQVN_N67, A2 => B1);
UQVB_B61 : AND4
	PORT MAP (Z0 => UQVN_N55, A0 => UQVN_N65, A1 => UQVN_N66, A2 => B0, 
	A3 => B2);
UQVB_B62 : OR7
	PORT MAP (Z0 => G012, A0 => UQVN_N52, A1 => UQVN_N51, A2 => UQVN_N50, 
	A3 => UQVN_N49, A4 => UQVN_N53, A5 => UQVN_N54, A6 => UQVN_N55);
UQVB_B63 : INV
	PORT MAP (ZN0 => UQVN_N68, A0 => B0);
UQVB_B64 : INV
	PORT MAP (ZN0 => UQVN_N66, A0 => A1);
UQVB_B65 : AND2
	PORT MAP (Z0 => UQVN_N46, A0 => A0, A1 => B1);
UQVB_B66 : AND2
	PORT MAP (Z0 => UQVN_N45, A0 => UQVN_N68, A1 => B1);
UQVB_B67 : OR3
	PORT MAP (Z0 => UQVN_N48, A0 => UQVN_N46, A1 => UQVN_N45, A2 => UQVN_N47);
UQVB_B68 : INV
	PORT MAP (ZN0 => UQVN_N70, A0 => B2);
UQVB_B69 : XOR2
	PORT MAP (Z0 => Z0, A0 => A0, A1 => B0);
UQVB_B70 : INV
	PORT MAP (ZN0 => UQVN_N67, A0 => A2);
UQVB_B71 : LXOR2
	PORT MAP (Z0 => Z2, A0 => A2, A1 => UQVN_N60);
UQVB_B72 : AND4
	PORT MAP (Z0 => UQVN_N59, A0 => UQVN_N65, A1 => B0, A2 => B1, 
	A3 => UQVN_N70);
UQVB_B73 : AND3
	PORT MAP (Z0 => UQVN_N58, A0 => A1, A1 => UQVN_N69, A2 => B2);
UQVB_B74 : AND4
	PORT MAP (Z0 => UQVN_N57, A0 => UQVN_N65, A1 => UQVN_N66, A2 => B0, 
	A3 => UQVN_N70);
UQVB_B75 : AND3
	PORT MAP (Z0 => UQVN_N56, A0 => UQVN_N68, A1 => UQVN_N69, A2 => B2);
UQVB_B76 : AND3
	PORT MAP (Z0 => UQVN_N64, A0 => A0, A1 => A1, A2 => B2);
UQVB_B77 : AND3
	PORT MAP (Z0 => UQVN_N63, A0 => A1, A1 => UQVN_N68, A2 => B2);
UQVB_B78 : AND3
	PORT MAP (Z0 => UQVN_N62, A0 => UQVN_N66, A1 => B1, A2 => UQVN_N70);
UQVB_B79 : AND3
	PORT MAP (Z0 => UQVN_N61, A0 => A0, A1 => UQVN_N69, A2 => B2);
UQVB_B80 : OR8
	PORT MAP (Z0 => UQVN_N60, A0 => UQVN_N64, A1 => UQVN_N63, A2 => UQVN_N62, 
	A3 => UQVN_N61, A4 => UQVN_N59, A5 => UQVN_N58, A6 => UQVN_N57, 
	A7 => UQVN_N56);
UQVB_B81 : INV
	PORT MAP (ZN0 => UQVN_N92, A0 => UQVN_N93);
UQVB_B82 : AND3
	PORT MAP (Z0 => UQVN_N73, A0 => UQVN_N93, A1 => UQVN_N89, A2 => UQVN_N88);
UQVB_B83 : AND3
	PORT MAP (Z0 => UQVN_N72, A0 => UQVN_N93, A1 => UQVN_N89, A2 => B6);
UQVB_B84 : AND3
	PORT MAP (Z0 => UQVN_N71, A0 => UQVN_N93, A1 => UQVN_N88, A2 => B7);
UQVB_B85 : AND3
	PORT MAP (Z0 => UQVN_N74, A0 => UQVN_N93, A1 => B7, A2 => B6);
UQVB_B86 : AND3
	PORT MAP (Z0 => UQVN_N75, A0 => UQVN_N89, A1 => UQVN_N88, A2 => B6);
UQVB_B87 : AND3
	PORT MAP (Z0 => UQVN_N77, A0 => UQVN_N88, A1 => B7, A2 => B6);
UQVB_B88 : AND2
	PORT MAP (Z0 => UQVN_N76, A0 => UQVN_N89, A1 => B7);
UQVB_B89 : OR7
	PORT MAP (Z0 => BO, A0 => UQVN_N73, A1 => UQVN_N72, A2 => UQVN_N71, 
	A3 => UQVN_N74, A4 => UQVN_N75, A5 => UQVN_N77, A6 => UQVN_N76);
UQVB_B90 : AND3
	PORT MAP (Z0 => UQVN_N78, A0 => A6, A1 => B7, A2 => UQVN_N92);
UQVB_B91 : AND3
	PORT MAP (Z0 => UQVN_N79, A0 => B7, A1 => UQVN_N90, A2 => UQVN_N92);
UQVB_B92 : AND3
	PORT MAP (Z0 => UQVN_N80, A0 => UQVN_N88, A1 => UQVN_N91, A2 => UQVN_N93);
UQVB_B93 : AND3
	PORT MAP (Z0 => UQVN_N81, A0 => UQVN_N91, A1 => B6, A2 => UQVN_N93);
UQVB_B94 : AND3
	PORT MAP (Z0 => UQVN_N82, A0 => A6, A1 => B7, A2 => UQVN_N90);
UQVB_B95 : AND3
	PORT MAP (Z0 => UQVN_N83, A0 => UQVN_N88, A1 => UQVN_N91, A2 => B6);
UQVB_B96 : OR6
	PORT MAP (Z0 => UQVN_N84, A0 => UQVN_N78, A1 => UQVN_N79, A2 => UQVN_N80, 
	A3 => UQVN_N81, A4 => UQVN_N82, A5 => UQVN_N83);
UQVB_B97 : LXOR2
	PORT MAP (Z0 => Z7, A0 => A7, A1 => UQVN_N84);
UQVB_B98 : INV
	PORT MAP (ZN0 => UQVN_N90, A0 => B6);
UQVB_B99 : INV
	PORT MAP (ZN0 => UQVN_N91, A0 => B7);
UQVB_B100 : INV
	PORT MAP (ZN0 => UQVN_N89, A0 => A7);
UQVB_B101 : INV
	PORT MAP (ZN0 => UQVN_N88, A0 => A6);
UQVB_B102 : XOR2
	PORT MAP (Z0 => Z6, A0 => A6, A1 => UQVN_N85);
UQVB_B103 : OR2
	PORT MAP (Z0 => UQVN_N85, A0 => UQVN_N86, A1 => UQVN_N87);
UQVB_B104 : AND2
	PORT MAP (Z0 => UQVN_N86, A0 => UQVN_N90, A1 => UQVN_N93);
UQVB_B105 : AND2
	PORT MAP (Z0 => UQVN_N87, A0 => UQVN_N92, A1 => B6);
END lattice_arch;
--*************************************************************
--*  Following Macros are used for 8K device                *--
--***********************************************************--

Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIID11E is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIID11E;

architecture LATTICE_ARCH of BIID11E is
    signal v107: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);
    
begin
    v110: XBIDI1
        port map(Z0 => v107,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    v111: XDFF1E
        port map(Q0 => Q0,
                 D0 => v107,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIID14E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIID14E;

architecture LATTICE_ARCH of BIID14E is
    signal v107, v117, v127, v137: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => v107, XB0 => XB0, A0 => A0, OE => OE);
    vv101: XBIDI1 port map(Z0 => v117, XB0 => XB1, A0 => A1, OE => OE);
    vv102: XBIDI1 port map(Z0 => v127, XB0 => XB2, A0 => A2, OE => OE);
    vv103: XBIDI1 port map(Z0 => v137, XB0 => XB3, A0 => A3, OE => OE);

    vv110: XDFF1E port map(Q0 => Q0, D0 => v107, CLK => CLK, EN => EN);
    vv111: XDFF1E port map(Q0 => Q1, D0 => v117, CLK => CLK, EN => EN);
    vv112: XDFF1E port map(Q0 => Q2, D0 => v127, CLK => CLK, EN => EN);
    vv113: XDFF1E port map(Q0 => Q3, D0 => v137, CLK => CLK, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIID91 is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic;
         CD: IN std_logic);
end BIID91;

architecture LATTICE_ARCH of BIID91 is
    signal v104: std_logic;
    
    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v107: XDFF2
        port map(Q0 => Q0,
                 D0 => v104,
                 CLK => CLK,
                 CD => CD);
    
    v108: XBIDI1
        port map(Z0 => v104,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIID91E is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic;
         CD: IN std_logic);
end BIID91E;

architecture LATTICE_ARCH of BIID91E is
    signal v108: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);
    
begin
    v111: XBIDI1
        port map(Z0 => v108,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    v112: XDFF2E
        port map(Q0 => Q0,
                 D0 => v108,
                 CLK => CLK,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIID94 is
    port(CD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIID94;

architecture LATTICE_ARCH of BIID94 is
    signal v104, v114, v124, v134: std_logic;

    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    vv100: XDFF2 port map(Q0 => Q0, D0 => v104, CLK => CLK, CD => CD);
    vv101: XDFF2 port map(Q0 => Q1, D0 => v114, CLK => CLK, CD => CD);
    vv102: XDFF2 port map(Q0 => Q2, D0 => v124, CLK => CLK, CD => CD);
    vv103: XDFF2 port map(Q0 => Q3, D0 => v134, CLK => CLK, CD => CD);

    vv110: XBIDI1 port map(Z0 => v104, XB0 => XB0, A0 => A0, OE => OE);
    vv111: XBIDI1 port map(Z0 => v114, XB0 => XB1, A0 => A1, OE => OE);
    vv112: XBIDI1 port map(Z0 => v124, XB0 => XB2, A0 => A2, OE => OE);
    vv113: XBIDI1 port map(Z0 => v134, XB0 => XB3, A0 => A3, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIID94E is
    port(CD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIID94E;

architecture LATTICE_ARCH of BIID94E is
    signal v108, v118, v128, v138: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => v108, XB0 => XB0, A0 => A0, OE => OE);
    vv101: XBIDI1 port map(Z0 => v118, XB0 => XB1, A0 => A1, OE => OE);
    vv102: XBIDI1 port map(Z0 => v128, XB0 => XB2, A0 => A2, OE => OE);
    vv103: XBIDI1 port map(Z0 => v138, XB0 => XB3, A0 => A3, OE => OE);

    vv110: XDFF2E port map(Q0 => Q0, D0 => v108, CLK => CLK, CD => CD, EN => EN);
    vv111: XDFF2E port map(Q0 => Q1, D0 => v118, CLK => CLK, CD => CD, EN => EN);
    vv112: XDFF2E port map(Q0 => Q2, D0 => v128, CLK => CLK, CD => CD, EN => EN);
    vv113: XDFF2E port map(Q0 => Q3, D0 => v138, CLK => CLK, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDA1 is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         OE: IN std_logic);
end BIIDA1;

architecture LATTICE_ARCH of BIIDA1 is
    signal v104: std_logic;
    
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v107: XDFF3
        port map(Q0 => Q0,
                 D0 => v104,
                 CLK => CLK,
                 SD => SD);
    
    v108: XBIDI1
        port map(Z0 => v104,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDA1E is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic;
         SD: IN std_logic);
end BIIDA1E;

architecture LATTICE_ARCH of BIIDA1E is
    signal v108: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);
    
begin
    v111: XBIDI1
        port map(Z0 => v108,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    v112: XDFF3E
        port map(Q0 => Q0,
                 D0 => v108,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDA4 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIIDA4;

architecture LATTICE_ARCH of BIIDA4 is
    signal v104, v114, v124, v134: std_logic;

    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    vv100: XDFF3 port map(Q0 => Q0, D0 => v104, CLK => CLK, SD => SD);
    vv101: XDFF3 port map(Q0 => Q1, D0 => v114, CLK => CLK, SD => SD);
    vv102: XDFF3 port map(Q0 => Q2, D0 => v124, CLK => CLK, SD => SD);
    vv103: XDFF3 port map(Q0 => Q3, D0 => v134, CLK => CLK, SD => SD);

    vv110: XBIDI1 port map(Z0 => v104, XB0 => XB0, A0 => A0, OE => OE);
    vv111: XBIDI1 port map(Z0 => v114, XB0 => XB1, A0 => A1, OE => OE);
    vv112: XBIDI1 port map(Z0 => v124, XB0 => XB2, A0 => A2, OE => OE);
    vv113: XBIDI1 port map(Z0 => v134, XB0 => XB3, A0 => A3, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDA4E is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIIDA4E;

architecture LATTICE_ARCH of BIIDA4E is
    signal v108, v118, v128, v138: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => v108, XB0 => XB0, A0 => A0, OE => OE);
    vv101: XBIDI1 port map(Z0 => v118, XB0 => XB1, A0 => A1, OE => OE);
    vv102: XBIDI1 port map(Z0 => v128, XB0 => XB2, A0 => A2, OE => OE);
    vv103: XBIDI1 port map(Z0 => v138, XB0 => XB3, A0 => A3, OE => OE);

    vv110: XDFF3E port map(Q0 => Q0, D0 => v108, CLK => CLK, SD => SD, EN => EN);
    vv111: XDFF3E port map(Q0 => Q1, D0 => v118, CLK => CLK, SD => SD, EN => EN);
    vv112: XDFF3E port map(Q0 => Q2, D0 => v128, CLK => CLK, SD => SD, EN => EN);
    vv113: XDFF3E port map(Q0 => Q3, D0 => v138, CLK => CLK, SD => SD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDB1 is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end BIIDB1;

architecture LATTICE_ARCH of BIIDB1 is
    signal v101: std_logic;
    
    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v104: XDFF4
        port map(Q0 => Q0,
                 D0 => v101,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v105: XBIDI1
        port map(Z0 => v101,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDB1E is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end BIIDB1E;

architecture LATTICE_ARCH of BIIDB1E is
    signal v105: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);
    
begin
    v108: XBIDI1
        port map(Z0 => v105,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    v109: XDFF4E
        port map(Q0 => Q0,
                 D0 => v105,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDB4 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIIDB4;

architecture LATTICE_ARCH of BIIDB4 is
    signal v101, v111, v121, v131: std_logic;

    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
   
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    vv100: XDFF4 port map(Q0 => Q0, D0 => v101, CLK => CLK, SD => SD, CD => CD);
    vv101: XDFF4 port map(Q0 => Q1, D0 => v111, CLK => CLK, SD => SD, CD => CD);
    vv102: XDFF4 port map(Q0 => Q2, D0 => v121, CLK => CLK, SD => SD, CD => CD);
    vv103: XDFF4 port map(Q0 => Q3, D0 => v131, CLK => CLK, SD => SD, CD => CD);

    vv110: XBIDI1 port map(Z0 => v101, XB0 => XB0, A0 => A0, OE => OE);
    vv111: XBIDI1 port map(Z0 => v111, XB0 => XB1, A0 => A1, OE => OE);
    vv112: XBIDI1 port map(Z0 => v121, XB0 => XB2, A0 => A2, OE => OE);
    vv113: XBIDI1 port map(Z0 => v131, XB0 => XB3, A0 => A3, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIDB4E is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIIDB4E;

architecture LATTICE_ARCH of BIIDB4E is
    signal v105, v115, v125, v135: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => v105, XB0 => XB0, A0 => A0, OE => OE);
    vv101: XBIDI1 port map(Z0 => v115, XB0 => XB1, A0 => A1, OE => OE);
    vv102: XBIDI1 port map(Z0 => v125, XB0 => XB2, A0 => A2, OE => OE);
    vv103: XBIDI1 port map(Z0 => v135, XB0 => XB3, A0 => A3, OE => OE);

    vv110: XDFF4E port map(Q0 => Q0, D0 => v105, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv111: XDFF4E port map(Q0 => Q1, D0 => v115, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv112: XDFF4E port map(Q0 => Q2, D0 => v125, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv113: XDFF4E port map(Q0 => Q3, D0 => v135, CLK => CLK, SD => SD, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIL91 is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic;
         CD: IN std_logic);
end BIIL91;

architecture LATTICE_ARCH of BIIL91 is
    signal v104: std_logic;
    
    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v107: XDL2
        port map(Q0 => Q0,
                 D0 => v104,
                 G => G,
                 CD => CD);
    
    v108: XBIDI1
        port map(Z0 => v104,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIIL94 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic;
         CD: IN std_logic);
end BIIL94;

architecture LATTICE_ARCH of BIIL94 is
    signal v104, v114, v124, v134: std_logic;

    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    v100: XDL2 port map(Q0 => Q0, D0 => v104, G => G, CD => CD);
    v101: XDL2 port map(Q0 => Q1, D0 => v114, G => G, CD => CD);
    v102: XDL2 port map(Q0 => Q2, D0 => v124, G => G, CD => CD);
    v103: XDL2 port map(Q0 => Q3, D0 => v134, G => G, CD => CD);

    v110: XBIDI1 port map(Z0 => v104, XB0 => XB0, A0 => A0, OE => OE);
    v111: XBIDI1 port map(Z0 => v114, XB0 => XB1, A0 => A1, OE => OE);
    v112: XBIDI1 port map(Z0 => v124, XB0 => XB2, A0 => A2, OE => OE);
    v113: XBIDI1 port map(Z0 => v134, XB0 => XB3, A0 => A3, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIILA1 is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic;
         SD: IN std_logic);
end BIILA1;

architecture LATTICE_ARCH of BIILA1 is
    signal v104: std_logic;
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v107: XDL3
        port map(Q0 => Q0,
                 D0 => v104,
                 G => G,
                 SD => SD);
    
    v108: XBIDI1
        port map(Z0 => v104,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIILA4 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic;
         SD: IN std_logic);
end BIILA4;

architecture LATTICE_ARCH of BIILA4 is
    signal v104, v114, v124, v134 : std_logic;

        component XDL3
            port(Q0: OUT std_logic;
                 D0: IN std_logic;
                 G: IN std_logic;
                 SD: IN std_logic);
        end component;
        for all: XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);
  
        component XBIDI1
            port(Z0: OUT std_logic;
                 XB0: INOUT std_logic;
                 A0: IN std_logic;
                 OE: IN std_logic);
        end component;
        for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    v100: XDL3 port map(Q0 => Q0, D0 => v104, G => G, SD => SD);
    v101: XDL3 port map(Q0 => Q1, D0 => v114, G => G, SD => SD);
    v102: XDL3 port map(Q0 => Q2, D0 => v124, G => G, SD => SD);
    v103: XDL3 port map(Q0 => Q3, D0 => v134, G => G, SD => SD);

    v110: XBIDI1 port map(Z0 => v104, XB0 => XB0, A0 => A0, OE => OE);
    v111: XBIDI1 port map(Z0 => v114, XB0 => XB1, A0 => A1, OE => OE);
    v112: XBIDI1 port map(Z0 => v124, XB0 => XB2, A0 => A2, OE => OE);
    v113: XBIDI1 port map(Z0 => v134, XB0 => XB3, A0 => A3, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIILB1 is
    port(Q0: OUT std_logic;
         XB0: INOUT std_logic;
         A0: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic);
end BIILB1;

architecture LATTICE_ARCH of BIILB1 is
    signal v102: std_logic;
    
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v105: XDL4
        port map(Q0 => Q0,
                 D0 => v102,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v106: XBIDI1
        port map(Z0 => v102,
                 XB0 => XB0,
                 A0 => A0,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIILB4 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic);
end BIILB4;

architecture LATTICE_ARCH of BIILB4 is
    signal v102, v112, v122, v132: std_logic;

    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
      
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    vv100: XDL4 port map(Q0 => Q0, D0 => v102, G => G, SD => SD, CD => CD);
    vv101: XDL4 port map(Q0 => Q1, D0 => v112, G => G, SD => SD, CD => CD);
    vv102: XDL4 port map(Q0 => Q2, D0 => v122, G => G, SD => SD, CD => CD);
    vv103: XDL4 port map(Q0 => Q3, D0 => v132, G => G, SD => SD, CD => CD);

    vv110: XBIDI1 port map(Z0 => v102, XB0 => XB0, A0 => A0, OE => OE);
    vv111: XBIDI1 port map(Z0 => v112, XB0 => XB1, A0 => A1, OE => OE);
    vv112: XBIDI1 port map(Z0 => v122, XB0 => XB2, A0 => A2, OE => OE);
    vv113: XBIDI1 port map(Z0 => v132, XB0 => XB3, A0 => A3, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD11 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD11;

architecture LATTICE_ARCH of BIOD11 is
    signal v101: std_logic;
    
    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
begin
    v104: XDFF1
        port map(Q0 => v101,
                 D0 => D0,
                 CLK => CLK);
    
    v105: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v101,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD11E is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD11E;

architecture LATTICE_ARCH of BIOD11E is
    signal v107: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);
    
begin
    v110: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v107,
                 OE => OE);
    
    v111: XDFF1E
        port map(Q0 => v107,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD14 is
    port(Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD14;

architecture LATTICE_ARCH of BIOD14 is
    signal v101, v111, v121, v131: std_logic;

    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);

begin

    vv100: XDFF1 port map(Q0 => v101, D0 => D0, CLK => CLK);
    vv101: XDFF1 port map(Q0 => v111, D0 => D1, CLK => CLK);
    vv102: XDFF1 port map(Q0 => v121, D0 => D2, CLK => CLK);
    vv103: XDFF1 port map(Q0 => v131, D0 => D3, CLK => CLK);

    vv110: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v101, OE => OE);
    vv111: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v111, OE => OE);
    vv112: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v121, OE => OE);
    vv113: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v131, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD14E is
    port(Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIOD14E;

architecture LATTICE_ARCH of BIOD14E is
    signal v107, v117, v127, v137: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v107, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v117, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v127, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v137, OE => OE);

    v110: XDFF1E port map(Q0 => v107, D0 => D0, CLK => CLK, EN => EN);
    v111: XDFF1E port map(Q0 => v117, D0 => D1, CLK => CLK, EN => EN);
    v112: XDFF1E port map(Q0 => v127, D0 => D2, CLK => CLK, EN => EN);
    v113: XDFF1E port map(Q0 => v137, D0 => D3, CLK => CLK, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD21 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CD: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD21;

architecture LATTICE_ARCH of BIOD21 is
    signal v104: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);
    
begin
    v107: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v104,
                 OE => OE);
    
    v108: XDFF2
        port map(Q0 => v104,
                 D0 => D0,
                 CLK => CLK,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD21E is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD21E;

architecture LATTICE_ARCH of BIOD21E is
    signal v108: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);
    
begin
    v111: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v108,
                 OE => OE);
    
    v112: XDFF2E
        port map(Q0 => v108,
                 D0 => D0,
                 CLK => CLK,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD24 is
    port(CD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD24;

architecture LATTICE_ARCH of BIOD24 is
    signal v104, v114, v124, v134: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v104, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v114, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v124, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v134, OE => OE);

    v110: XDFF2 port map(Q0 => v104, D0 => D0, CLK => CLK, CD => CD);
    v111: XDFF2 port map(Q0 => v114, D0 => D1, CLK => CLK, CD => CD);
    v112: XDFF2 port map(Q0 => v124, D0 => D2, CLK => CLK, CD => CD);
    v113: XDFF2 port map(Q0 => v134, D0 => D3, CLK => CLK, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD24E is
    port(CD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIOD24E;

architecture LATTICE_ARCH of BIOD24E is
    signal v108, v118, v128, v138: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v108, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v118, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v128, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v138, OE => OE);

    v110: XDFF2E port map(Q0 => v108, D0 => D0, CLK => CLK, CD => CD, EN => EN);
    v111: XDFF2E port map(Q0 => v118, D0 => D1, CLK => CLK, CD => CD, EN => EN);
    v112: XDFF2E port map(Q0 => v128, D0 => D2, CLK => CLK, CD => CD, EN => EN);
    v113: XDFF2E port map(Q0 => v138, D0 => D3, CLK => CLK, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD31 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         SD: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD31;

architecture LATTICE_ARCH of BIOD31 is
    signal v104: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);
    
begin
    v107: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v104,
                 OE => OE);
    
    v108: XDFF3
        port map(Q0 => v104,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD31E is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD31E;

architecture LATTICE_ARCH of BIOD31E is
    signal v108: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);
    
begin
    v111: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v108,
                 OE => OE);
    
    v112: XDFF3E
        port map(Q0 => v108,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD34 is
    port(SD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD34;

architecture LATTICE_ARCH of BIOD34 is
    signal v104, v114, v124, v134: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v104, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v114, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v124, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v134, OE => OE);

    v110: XDFF3 port map(Q0 => v104, D0 => D0, CLK => CLK, SD => SD);
    v111: XDFF3 port map(Q0 => v114, D0 => D1, CLK => CLK, SD => SD);
    v112: XDFF3 port map(Q0 => v124, D0 => D2, CLK => CLK, SD => SD);
    v113: XDFF3 port map(Q0 => v134, D0 => D3, CLK => CLK, SD => SD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD34E is
    port(SD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIOD34E;

architecture LATTICE_ARCH of BIOD34E is
    signal v108, v118, v128, v138: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v108, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v118, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v128, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v138, OE => OE);

    v110: XDFF3E port map(Q0 => v108, D0 => D0, CLK => CLK, SD => SD, EN => EN);
    v111: XDFF3E port map(Q0 => v118, D0 => D1, CLK => CLK, SD => SD, EN => EN);
    v112: XDFF3E port map(Q0 => v128, D0 => D2, CLK => CLK, SD => SD, EN => EN);
    v113: XDFF3E port map(Q0 => v138, D0 => D3, CLK => CLK, SD => SD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD41 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD41;

architecture LATTICE_ARCH of BIOD41 is
    signal v101: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
    
begin
    v104: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v101,
                 OE => OE);
    
    v105: XDFF4
        port map(Q0 => v101,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD41E is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD41E;

architecture LATTICE_ARCH of BIOD41E is
    signal v105: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);
    
begin
    v108: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v105,
                 OE => OE);
    
    v109: XDFF4E
        port map(Q0 => v105,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD44 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end BIOD44;

architecture LATTICE_ARCH of BIOD44 is
    signal v101, v111, v121, v131: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v101, OE => OE);
    vv101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v111, OE => OE);
    vv102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v121, OE => OE);
    vv103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v131, OE => OE);

    vv110: XDFF4 port map(Q0 => v101, D0 => D0, CLK => CLK, SD => SD, CD => CD);
    vv111: XDFF4 port map(Q0 => v111, D0 => D1, CLK => CLK, SD => SD, CD => CD);
    vv112: XDFF4 port map(Q0 => v121, D0 => D2, CLK => CLK, SD => SD, CD => CD);
    vv113: XDFF4 port map(Q0 => v131, D0 => D3, CLK => CLK, SD => SD, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOD44E is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end BIOD44E;

architecture LATTICE_ARCH of BIOD44E is
    signal v105, v115, v125, v135: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v105, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v115, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v125, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v135, OE => OE);

    v110: XDFF4E port map(Q0 => v105, D0 => D0, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v111: XDFF4E port map(Q0 => v115, D0 => D1, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v112: XDFF4E port map(Q0 => v125, D0 => D2, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v113: XDFF4E port map(Q0 => v135, D0 => D3, CLK => CLK, SD => SD, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL11 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL11;

architecture LATTICE_ARCH of BIOL11 is
    signal v101: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);
    
begin
    v104: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v101,
                 OE => OE);
    
    v105: XDL1
        port map(Q0 => v101,
                 D0 => D0,
                 G => G);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL14 is
    port(Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL14;

architecture LATTICE_ARCH of BIOL14 is
    signal v101, v111, v121, v131 : std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v101, OE => OE);
    vv101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v111, OE => OE);
    vv102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v121, OE => OE);
    vv103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v131, OE => OE);

    vv110: XDL1 port map(Q0 => v101, D0 => D0, G => G);
    vv111: XDL1 port map(Q0 => v111, D0 => D1, G => G);
    vv112: XDL1 port map(Q0 => v121, D0 => D2, G => G);
    vv113: XDL1 port map(Q0 => v131, D0 => D3, G => G);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL21 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CD: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL21;

architecture LATTICE_ARCH of BIOL21 is
    signal v104: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);
    
begin
    v107: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v104,
                 OE => OE);
    
    v108: XDL2
        port map(Q0 => v104,
                 D0 => D0,
                 G => G,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL24 is
    port(CD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL24;

architecture LATTICE_ARCH of BIOL24 is
    signal v104, v114, v124, v134: std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
   
    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v104, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v114, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v124, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v134, OE => OE);

    v110: XDL2 port map(Q0 => v104, D0 => D0, G => G, CD => CD);
    v111: XDL2 port map(Q0 => v114, D0 => D1, G => G, CD => CD);
    v112: XDL2 port map(Q0 => v124, D0 => D2, G => G, CD => CD);
    v113: XDL2 port map(Q0 => v134, D0 => D3, G => G, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL31 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         SD: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL31;

architecture LATTICE_ARCH of BIOL31 is
    signal v104: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);
    
begin
    v107: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v104,
                 OE => OE);
    
    v108: XDL3
        port map(Q0 => v104,
                 D0 => D0,
                 G => G,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL34 is
    port(SD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL34;

architecture LATTICE_ARCH of BIOL34 is
    signal v104, v114, v124, v134 : std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);

begin

    v100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v104, OE => OE);
    v101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v114, OE => OE);
    v102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v124, OE => OE);
    v103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v134, OE => OE);

    v110: XDL3 port map(Q0 => v104, D0 => D0, G => G, SD => SD);
    v111: XDL3 port map(Q0 => v114, D0 => D1, G => G, SD => SD);
    v112: XDL3 port map(Q0 => v124, D0 => D2, G => G, SD => SD);
    v113: XDL3 port map(Q0 => v134, D0 => D3, G => G, SD => SD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL41 is
    port(Z0: OUT std_logic;
         XB0: INOUT std_logic;
         D0: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL41;

architecture LATTICE_ARCH of BIOL41 is
    signal v102: std_logic;
    
    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
    
begin
    v105: XBIDI1
        port map(Z0 => Z0,
                 XB0 => XB0,
                 A0 => v102,
                 OE => OE);
    
    v106: XDL4
        port map(Q0 => v102,
                 D0 => D0,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity BIOL44 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Z0: OUT std_logic;
         Z1: OUT std_logic;
         Z2: OUT std_logic;
         Z3: OUT std_logic;
         XB0: INOUT std_logic;
         XB1: INOUT std_logic;
         XB2: INOUT std_logic;
         XB3: INOUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end BIOL44;

architecture LATTICE_ARCH of BIOL44 is
    signal v102, v112, v122, v132 : std_logic;

    component XBIDI1
        port(Z0: OUT std_logic;
             XB0: INOUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XBIDI1 use entity LAT_VHD.XBIDI1(LATTICE_ARCH);
    
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);

begin

    vv100: XBIDI1 port map(Z0 => Z0, XB0 => XB0, A0 => v102, OE => OE);
    vv101: XBIDI1 port map(Z0 => Z1, XB0 => XB1, A0 => v112, OE => OE);
    vv102: XBIDI1 port map(Z0 => Z2, XB0 => XB2, A0 => v122, OE => OE);
    vv103: XBIDI1 port map(Z0 => Z3, XB0 => XB3, A0 => v132, OE => OE);

    vv110: XDL4 port map(Q0 => v102, D0 => D0, G => G, SD => SD, CD => CD);
    vv111: XDL4 port map(Q0 => v112, D0 => D1, G => G, SD => SD, CD => CD);
    vv112: XDL4 port map(Q0 => v122, D0 => D2, G => G, SD => SD, CD => CD);
    vv113: XDL4 port map(Q0 => v132, D0 => D3, G => G, SD => SD, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBD84 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic);
end CBD84;

architecture LATTICE_ARCH of CBD84 is
    signal QI: std_logic_vector(0 to 3);
    signal v115: std_logic_vector(0 to 3);
    signal v103: std_logic;
    signal v110: std_logic;
    signal v108: std_logic;
    signal v107: std_logic;
    signal v106: std_logic;
    signal v105: std_logic;
    signal v104: std_logic;
    signal v109: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v137: FDC1
        port map(Q0 => QI(0),
                 D0 => v107,
                 CLK => CLK,
                 SD => SD);
    
    v138: FDC1
        port map(Q0 => QI(1),
                 D0 => v108,
                 CLK => CLK,
                 SD => SD);
    
    v139: AND2
        port map(Z0 => v103,
                 A0 => CAI,
                 A1 => EN);
    
    v140: AND3
        port map(Z0 => v104,
                 A0 => v115(0),
                 A1 => CAI,
                 A2 => EN);
    
    v141: AND4
        port map(Z0 => v105,
                 A0 => v115(0),
                 A1 => v115(1),
                 A2 => CAI,
                 A3 => EN);
    
    v142: AND5
        port map(Z0 => v106,
                 A0 => v115(0),
                 A1 => v115(1),
                 A2 => v115(2),
                 A3 => CAI,
                 A4 => EN);
    
    v143: AND6
        port map(Z0 => CAO,
                 A0 => v115(0),
                 A1 => v115(1),
                 A2 => v115(2),
                 A3 => v115(3),
                 A4 => CAI,
                 A5 => EN);
    
    v144: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v145: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v146: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v147: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v148: INV
        port map(ZN0 => v115(0),
                 A0 => QI(0));
    
    v149: INV
        port map(ZN0 => v115(1),
                 A0 => QI(1));
    
    v150: INV
        port map(ZN0 => v115(2),
                 A0 => QI(2));
    
    v151: INV
        port map(ZN0 => v115(3),
                 A0 => QI(3));
    
    v152: FDC1
        port map(Q0 => QI(2),
                 D0 => v109,
                 CLK => CLK,
                 SD => SD);
    
    v153: FDC1
        port map(Q0 => QI(3),
                 D0 => v110,
                 CLK => CLK,
                 SD => SD);
    
    v154: LXOR2
        port map(Z0 => v107,
                 A0 => QI(0),
                 A1 => v103);
    
    v155: LXOR2
        port map(Z0 => v108,
                 A0 => QI(1),
                 A1 => v104);
    
    v156: LXOR2
        port map(Z0 => v109,
                 A0 => QI(2),
                 A1 => v105);
    
    v157: LXOR2
        port map(Z0 => v110,
                 A0 => QI(3),
                 A1 => v106);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBD88 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic);
end CBD88;

architecture LATTICE_ARCH of CBD88 is
    signal QI: std_logic_vector(0 to 7);
    signal v129: std_logic_vector(0 to 7);
    signal v105: std_logic;
    signal v119: std_logic;
    signal v116: std_logic;
    signal v114: std_logic;
    signal v111: std_logic;
    signal v113: std_logic;
    signal v108: std_logic;
    signal v107: std_logic;
    signal v106: std_logic;
    signal v117: std_logic;
    signal v115: std_logic;
    signal v120: std_logic;
    signal v112: std_logic;
    signal v109: std_logic;
    signal v118: std_logic;
    signal v110: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v171: FDC1
        port map(Q0 => QI(0),
                 D0 => v113,
                 CLK => CLK,
                 SD => SD);
    
    v172: FDC1
        port map(Q0 => QI(1),
                 D0 => v114,
                 CLK => CLK,
                 SD => SD);
    
    v173: AND10
        port map(Z0 => CAO,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v129(3),
                 A4 => v129(4),
                 A5 => v129(5),
                 A6 => v129(6),
                 A7 => v129(7),
                 A8 => CAI,
                 A9 => EN);
    
    v174: AND2
        port map(Z0 => v105,
                 A0 => CAI,
                 A1 => EN);
    
    v175: AND3
        port map(Z0 => v106,
                 A0 => v129(0),
                 A1 => CAI,
                 A2 => EN);
    
    v176: AND4
        port map(Z0 => v107,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => CAI,
                 A3 => EN);
    
    v177: AND5
        port map(Z0 => v108,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => CAI,
                 A4 => EN);
    
    v178: AND6
        port map(Z0 => v109,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v129(3),
                 A4 => CAI,
                 A5 => EN);
    
    v179: AND7
        port map(Z0 => v110,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v129(3),
                 A4 => v129(4),
                 A5 => CAI,
                 A6 => EN);
    
    v180: AND8
        port map(Z0 => v111,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v129(3),
                 A4 => v129(4),
                 A5 => v129(5),
                 A6 => CAI,
                 A7 => EN);
    
    v181: AND9
        port map(Z0 => v112,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v129(3),
                 A4 => v129(4),
                 A5 => v129(5),
                 A6 => v129(6),
                 A7 => CAI,
                 A8 => EN);
    
    v182: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v183: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v184: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v185: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v186: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v187: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v188: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v189: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v190: INV
        port map(ZN0 => v129(0),
                 A0 => QI(0));
    
    v191: INV
        port map(ZN0 => v129(1),
                 A0 => QI(1));
    
    v192: INV
        port map(ZN0 => v129(2),
                 A0 => QI(2));
    
    v193: INV
        port map(ZN0 => v129(3),
                 A0 => QI(3));
    
    v194: INV
        port map(ZN0 => v129(4),
                 A0 => QI(4));
    
    v195: INV
        port map(ZN0 => v129(5),
                 A0 => QI(5));
    
    v196: INV
        port map(ZN0 => v129(6),
                 A0 => QI(6));
    
    v197: INV
        port map(ZN0 => v129(7),
                 A0 => QI(7));
    
    v198: FDC1
        port map(Q0 => QI(2),
                 D0 => v115,
                 CLK => CLK,
                 SD => SD);
    
    v199: FDC1
        port map(Q0 => QI(3),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD);
    
    v200: LXOR2
        port map(Z0 => v113,
                 A0 => QI(0),
                 A1 => v105);
    
    v201: LXOR2
        port map(Z0 => v114,
                 A0 => QI(1),
                 A1 => v106);
    
    v202: LXOR2
        port map(Z0 => v115,
                 A0 => QI(2),
                 A1 => v107);
    
    v203: LXOR2
        port map(Z0 => v116,
                 A0 => QI(3),
                 A1 => v108);
    
    v204: LXOR2
        port map(Z0 => v117,
                 A0 => QI(4),
                 A1 => v109);
    
    v205: FDC1
        port map(Q0 => QI(4),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD);
    
    v206: LXOR2
        port map(Z0 => v118,
                 A0 => QI(5),
                 A1 => v110);
    
    v207: FDC1
        port map(Q0 => QI(5),
                 D0 => v118,
                 CLK => CLK,
                 SD => SD);
    
    v208: FDC1
        port map(Q0 => QI(6),
                 D0 => v119,
                 CLK => CLK,
                 SD => SD);
    
    v209: LXOR2
        port map(Z0 => v119,
                 A0 => QI(6),
                 A1 => v111);
    
    v210: LXOR2
        port map(Z0 => v120,
                 A0 => QI(7),
                 A1 => v112);
    
    v211: FDC1
        port map(Q0 => QI(7),
                 D0 => v120,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBD94 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBD94;

architecture LATTICE_ARCH of CBD94 is
    signal QI: std_logic_vector(0 to 3);
    signal v112: std_logic_vector(0 to 3);
    signal v100: std_logic;
    signal v107: std_logic;
    signal v105: std_logic;
    signal v104: std_logic;
    signal v103: std_logic;
    signal v102: std_logic;
    signal v101: std_logic;
    signal v106: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v134: FDE1
        port map(Q0 => QI(0),
                 D0 => v104,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v135: FDE1
        port map(Q0 => QI(1),
                 D0 => v105,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v136: AND2
        port map(Z0 => v100,
                 A0 => CAI,
                 A1 => EN);
    
    v137: AND3
        port map(Z0 => v101,
                 A0 => v112(0),
                 A1 => CAI,
                 A2 => EN);
    
    v138: AND4
        port map(Z0 => v102,
                 A0 => v112(0),
                 A1 => v112(1),
                 A2 => CAI,
                 A3 => EN);
    
    v139: AND5
        port map(Z0 => v103,
                 A0 => v112(0),
                 A1 => v112(1),
                 A2 => v112(2),
                 A3 => CAI,
                 A4 => EN);
    
    v140: AND6
        port map(Z0 => CAO,
                 A0 => v112(0),
                 A1 => v112(1),
                 A2 => v112(2),
                 A3 => v112(3),
                 A4 => CAI,
                 A5 => EN);
    
    v141: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v142: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v143: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v144: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v145: INV
        port map(ZN0 => v112(0),
                 A0 => QI(0));
    
    v146: INV
        port map(ZN0 => v112(1),
                 A0 => QI(1));
    
    v147: INV
        port map(ZN0 => v112(2),
                 A0 => QI(2));
    
    v148: INV
        port map(ZN0 => v112(3),
                 A0 => QI(3));
    
    v149: FDE1
        port map(Q0 => QI(2),
                 D0 => v106,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v150: FDE1
        port map(Q0 => QI(3),
                 D0 => v107,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v151: LXOR2
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => v100);
    
    v152: LXOR2
        port map(Z0 => v105,
                 A0 => QI(1),
                 A1 => v101);
    
    v153: LXOR2
        port map(Z0 => v106,
                 A0 => QI(2),
                 A1 => v102);
    
    v154: LXOR2
        port map(Z0 => v107,
                 A0 => QI(3),
                 A1 => v103);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBD98 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBD98;

architecture LATTICE_ARCH of CBD98 is
    signal QI: std_logic_vector(0 to 7);
    signal v126: std_logic_vector(0 to 7);
    signal v102: std_logic;
    signal v116: std_logic;
    signal v113: std_logic;
    signal v111: std_logic;
    signal v108: std_logic;
    signal v110: std_logic;
    signal v105: std_logic;
    signal v104: std_logic;
    signal v103: std_logic;
    signal v114: std_logic;
    signal v112: std_logic;
    signal v117: std_logic;
    signal v109: std_logic;
    signal v106: std_logic;
    signal v115: std_logic;
    signal v107: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v168: FDE1
        port map(Q0 => QI(0),
                 D0 => v110,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v169: FDE1
        port map(Q0 => QI(1),
                 D0 => v111,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v170: AND10
        port map(Z0 => CAO,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => v126(2),
                 A3 => v126(3),
                 A4 => v126(4),
                 A5 => v126(5),
                 A6 => v126(6),
                 A7 => v126(7),
                 A8 => CAI,
                 A9 => EN);
    
    v171: AND2
        port map(Z0 => v102,
                 A0 => CAI,
                 A1 => EN);
    
    v172: AND3
        port map(Z0 => v103,
                 A0 => v126(0),
                 A1 => CAI,
                 A2 => EN);
    
    v173: AND4
        port map(Z0 => v104,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => CAI,
                 A3 => EN);
    
    v174: AND5
        port map(Z0 => v105,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => v126(2),
                 A3 => CAI,
                 A4 => EN);
    
    v175: AND6
        port map(Z0 => v106,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => v126(2),
                 A3 => v126(3),
                 A4 => CAI,
                 A5 => EN);
    
    v176: AND7
        port map(Z0 => v107,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => v126(2),
                 A3 => v126(3),
                 A4 => v126(4),
                 A5 => CAI,
                 A6 => EN);
    
    v177: AND8
        port map(Z0 => v108,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => v126(2),
                 A3 => v126(3),
                 A4 => v126(4),
                 A5 => v126(5),
                 A6 => CAI,
                 A7 => EN);
    
    v178: AND9
        port map(Z0 => v109,
                 A0 => v126(0),
                 A1 => v126(1),
                 A2 => v126(2),
                 A3 => v126(3),
                 A4 => v126(4),
                 A5 => v126(5),
                 A6 => v126(6),
                 A7 => CAI,
                 A8 => EN);
    
    v179: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v180: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v181: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v182: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v183: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v184: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v185: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v186: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v187: INV
        port map(ZN0 => v126(0),
                 A0 => QI(0));
    
    v188: INV
        port map(ZN0 => v126(1),
                 A0 => QI(1));
    
    v189: INV
        port map(ZN0 => v126(2),
                 A0 => QI(2));
    
    v190: INV
        port map(ZN0 => v126(3),
                 A0 => QI(3));
    
    v191: INV
        port map(ZN0 => v126(4),
                 A0 => QI(4));
    
    v192: INV
        port map(ZN0 => v126(5),
                 A0 => QI(5));
    
    v193: INV
        port map(ZN0 => v126(6),
                 A0 => QI(6));
    
    v194: INV
        port map(ZN0 => v126(7),
                 A0 => QI(7));
    
    v195: FDE1
        port map(Q0 => QI(2),
                 D0 => v112,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v196: FDE1
        port map(Q0 => QI(3),
                 D0 => v113,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v197: LXOR2
        port map(Z0 => v110,
                 A0 => QI(0),
                 A1 => v102);
    
    v198: LXOR2
        port map(Z0 => v111,
                 A0 => QI(1),
                 A1 => v103);
    
    v199: LXOR2
        port map(Z0 => v112,
                 A0 => QI(2),
                 A1 => v104);
    
    v200: LXOR2
        port map(Z0 => v113,
                 A0 => QI(3),
                 A1 => v105);
    
    v201: LXOR2
        port map(Z0 => v114,
                 A0 => QI(4),
                 A1 => v106);
    
    v202: FDE1
        port map(Q0 => QI(4),
                 D0 => v114,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v203: LXOR2
        port map(Z0 => v115,
                 A0 => QI(5),
                 A1 => v107);
    
    v204: FDE1
        port map(Q0 => QI(5),
                 D0 => v115,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v205: FDE1
        port map(Q0 => QI(6),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v206: LXOR2
        port map(Z0 => v116,
                 A0 => QI(6),
                 A1 => v108);
    
    v207: LXOR2
        port map(Z0 => v117,
                 A0 => QI(7),
                 A1 => v109);
    
    v208: FDE1
        port map(Q0 => QI(7),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBDA16 is
    port(CAI: IN std_logic;
         CAO: OUT std_logic;
         CD: IN std_logic;
         CLK: IN std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D10: IN std_logic;
         D11: IN std_logic;
         D12: IN std_logic;
         D13: IN std_logic;
         D14: IN std_logic;
         D15: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         D8: IN std_logic;
         D9: IN std_logic;
         EN: IN std_logic;
         LD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q10: OUT std_logic;
         Q11: OUT std_logic;
         Q12: OUT std_logic;
         Q13: OUT std_logic;
         Q14: OUT std_logic;
         Q15: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         Q8: OUT std_logic;
         Q9: OUT std_logic;
         SD: IN std_logic);
end CBDA16;

architecture LATTICE_ARCH of CBDA16 is
    signal QI: std_logic_vector(0 to 15);
    signal v205: std_logic_vector(0 to 15);
    signal v125: std_logic;
    signal v113: std_logic;
    signal v136: std_logic;
    signal v111: std_logic;
    signal v152: std_logic;
    signal v133: std_logic;
    signal v121: std_logic;
    signal v143: std_logic;
    signal v135: std_logic;
    signal v120: std_logic;
    signal v112: std_logic;
    signal v179: std_logic;
    signal v159: std_logic;
    signal v122: std_logic;
    signal v129: std_logic;
    signal v127: std_logic;
    signal v114: std_logic;
    signal v183: std_logic;
    signal v146: std_logic;
    signal v126: std_logic;
    signal v124: std_logic;
    signal v162: std_logic;
    signal v150: std_logic;
    signal v134: std_logic;
    signal v123: std_logic;
    signal v119: std_logic;
    signal v116: std_logic;
    signal v166: std_logic;
    signal v131: std_logic;
    signal v128: std_logic;
    signal v115: std_logic;
    signal v186: std_logic;
    signal v167: std_logic;
    signal v132: std_logic;
    signal v188: std_logic;
    signal v117: std_logic;
    signal v118: std_logic;
    signal v110: std_logic;
    signal v104: std_logic;
    signal v130: std_logic;
    signal v151: std_logic;
    signal v139: std_logic;
    signal v178: std_logic;
    signal v155: std_logic;
    signal v140: std_logic;
    signal v156: std_logic;
    signal v181: std_logic;
    signal v173: std_logic;
    signal v105: std_logic;
    signal v182: std_logic;
    signal v147: std_logic;
    signal v106: std_logic;
    signal v163: std_logic;
    signal v141: std_logic;
    signal v107: std_logic;
    signal v157: std_logic;
    signal v148: std_logic;
    signal v142: std_logic;
    signal v108: std_logic;
    signal v187: std_logic;
    signal v169: std_logic;
    signal v164: std_logic;
    signal v158: std_logic;
    signal v144: std_logic;
    signal v137: std_logic;
    signal v174: std_logic;
    signal v170: std_logic;
    signal v160: std_logic;
    signal v153: std_logic;
    signal v149: std_logic;
    signal v138: std_logic;
    signal v109: std_logic;
    signal v168: std_logic;
    signal v165: std_logic;
    signal v154: std_logic;
    signal v184: std_logic;
    signal v175: std_logic;
    signal v171: std_logic;
    signal v180: std_logic;
    signal v172: std_logic;
    signal v145: std_logic;
    signal v176: std_logic;
    signal v161: std_logic;
    signal v185: std_logic;
    signal v177: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND18
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic;
             A15: IN std_logic;
             A16: IN std_logic;
             A17: IN std_logic);
    end component;
    for all : AND18 use entity LAT_VHD.AND18(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND11
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic);
    end component;
    for all : AND11 use entity LAT_VHD.AND11(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component AND12
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic);
    end component;
    for all : AND12 use entity LAT_VHD.AND12(LATTICE_ARCH);
    
    component AND13
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic);
    end component;
    for all : AND13 use entity LAT_VHD.AND13(LATTICE_ARCH);
    
    component AND14
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic);
    end component;
    for all : AND14 use entity LAT_VHD.AND14(LATTICE_ARCH);
    
    component AND15
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic);
    end component;
    for all : AND15 use entity LAT_VHD.AND15(LATTICE_ARCH);
    
    component AND16
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic;
             A15: IN std_logic);
    end component;
    for all : AND16 use entity LAT_VHD.AND16(LATTICE_ARCH);
    
    component AND17
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic;
             A15: IN std_logic;
             A16: IN std_logic);
    end component;
    for all : AND17 use entity LAT_VHD.AND17(LATTICE_ARCH);
    
begin
    v340: FDE1
        port map(Q0 => QI(0),
                 D0 => v126,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v341: FDE1
        port map(Q0 => QI(1),
                 D0 => v127,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v342: AND2
        port map(Z0 => v111,
                 A0 => D0,
                 A1 => LD);
    
    v343: AND3
        port map(Z0 => v112,
                 A0 => v125,
                 A1 => CAI,
                 A2 => EN);
    
    v344: AND2
        port map(Z0 => v114,
                 A0 => D1,
                 A1 => LD);
    
    v345: AND2
        port map(Z0 => v117,
                 A0 => D2,
                 A1 => LD);
    
    v346: AND2
        port map(Z0 => v121,
                 A0 => D3,
                 A1 => LD);
    
    v347: AND4
        port map(Z0 => v105,
                 A0 => v205(0),
                 A1 => CAI,
                 A2 => v125,
                 A3 => EN);
    
    v348: AND5
        port map(Z0 => v120,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v125,
                 A3 => CAI,
                 A4 => EN);
    
    v349: AND6
        port map(Z0 => v124,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v125,
                 A4 => CAI,
                 A5 => EN);
    
    v350: AND18
        port map(Z0 => CAO,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v205(10),
                 A11 => v205(11),
                 A12 => v205(12),
                 A13 => v205(13),
                 A14 => v205(14),
                 A15 => v205(15),
                 A16 => CAI,
                 A17 => EN);
    
    v351: AND2
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => v125);
    
    v352: OR2
        port map(Z0 => v113,
                 A0 => v111,
                 A1 => v112);
    
    v353: BUF
        port map(Z0 => Q15,
                 A0 => QI(15));
    
    v354: BUF
        port map(Z0 => Q11,
                 A0 => QI(11));
    
    v355: BUF
        port map(Z0 => Q9,
                 A0 => QI(9));
    
    v356: BUF
        port map(Z0 => Q8,
                 A0 => QI(8));
    
    v357: BUF
        port map(Z0 => Q14,
                 A0 => QI(14));
    
    v358: BUF
        port map(Z0 => Q13,
                 A0 => QI(13));
    
    v359: BUF
        port map(Z0 => Q12,
                 A0 => QI(12));
    
    v360: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v361: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v362: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v363: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v364: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v365: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v366: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v367: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v368: BUF
        port map(Z0 => Q10,
                 A0 => QI(10));
    
    v369: AND2
        port map(Z0 => v115,
                 A0 => QI(1),
                 A1 => v125);
    
    v370: OR2
        port map(Z0 => v116,
                 A0 => v114,
                 A1 => v105);
    
    v371: AND2
        port map(Z0 => v118,
                 A0 => QI(2),
                 A1 => v125);
    
    v372: OR2
        port map(Z0 => v119,
                 A0 => v117,
                 A1 => v120);
    
    v373: AND2
        port map(Z0 => v122,
                 A0 => QI(3),
                 A1 => v125);
    
    v374: OR2
        port map(Z0 => v123,
                 A0 => v121,
                 A1 => v124);
    
    v375: OR2
        port map(Z0 => v110,
                 A0 => v106,
                 A1 => v108);
    
    v376: AND2
        port map(Z0 => v109,
                 A0 => QI(4),
                 A1 => v125);
    
    v377: LXOR2
        port map(Z0 => v107,
                 A0 => v109,
                 A1 => v110);
    
    v378: FDE1
        port map(Q0 => QI(4),
                 D0 => v107,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v379: AND2
        port map(Z0 => v106,
                 A0 => D4,
                 A1 => LD);
    
    v380: AND7
        port map(Z0 => v108,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v125,
                 A5 => CAI,
                 A6 => EN);
    
    v381: INV
        port map(ZN0 => v205(0),
                 A0 => QI(0));
    
    v382: INV
        port map(ZN0 => v205(1),
                 A0 => QI(1));
    
    v383: INV
        port map(ZN0 => v205(2),
                 A0 => QI(2));
    
    v384: INV
        port map(ZN0 => v205(3),
                 A0 => QI(3));
    
    v385: INV
        port map(ZN0 => v205(4),
                 A0 => QI(4));
    
    v386: FDE1
        port map(Q0 => QI(2),
                 D0 => v128,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v387: FDE1
        port map(Q0 => QI(3),
                 D0 => v129,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v388: LXOR2
        port map(Z0 => v126,
                 A0 => v104,
                 A1 => v113);
    
    v389: LXOR2
        port map(Z0 => v127,
                 A0 => v115,
                 A1 => v116);
    
    v390: INV
        port map(ZN0 => v125,
                 A0 => LD);
    
    v391: LXOR2
        port map(Z0 => v128,
                 A0 => v118,
                 A1 => v119);
    
    v392: LXOR2
        port map(Z0 => v129,
                 A0 => v122,
                 A1 => v123);
    
    v393: AND10
        port map(Z0 => v136,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v143,
                 A8 => CAI,
                 A9 => EN);
    
    v394: INV
        port map(ZN0 => v143,
                 A0 => LD);
    
    v395: AND2
        port map(Z0 => v141,
                 A0 => QI(5),
                 A1 => v143);
    
    v396: OR2
        port map(Z0 => v148,
                 A0 => v137,
                 A1 => v149);
    
    v397: AND2
        port map(Z0 => v150,
                 A0 => QI(6),
                 A1 => v143);
    
    v398: OR2
        port map(Z0 => v145,
                 A0 => v130,
                 A1 => v147);
    
    v399: AND2
        port map(Z0 => v138,
                 A0 => QI(7),
                 A1 => v143);
    
    v400: OR2
        port map(Z0 => v144,
                 A0 => v140,
                 A1 => v136);
    
    v401: OR2
        port map(Z0 => v134,
                 A0 => v131,
                 A1 => v135);
    
    v402: AND2
        port map(Z0 => v133,
                 A0 => QI(8),
                 A1 => v143);
    
    v403: LXOR2
        port map(Z0 => v132,
                 A0 => v133,
                 A1 => v134);
    
    v404: AND2
        port map(Z0 => v131,
                 A0 => D8,
                 A1 => LD);
    
    v405: FDE1
        port map(Q0 => QI(8),
                 D0 => v132,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v406: AND11
        port map(Z0 => v135,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v143,
                 A9 => CAI,
                 A10 => EN);
    
    v407: INV
        port map(ZN0 => v205(5),
                 A0 => QI(5));
    
    v408: INV
        port map(ZN0 => v205(6),
                 A0 => QI(6));
    
    v409: INV
        port map(ZN0 => v205(7),
                 A0 => QI(7));
    
    v410: INV
        port map(ZN0 => v205(8),
                 A0 => QI(8));
    
    v411: AND8
        port map(Z0 => v149,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v143,
                 A6 => CAI,
                 A7 => EN);
    
    v412: AND2
        port map(Z0 => v137,
                 A0 => D5,
                 A1 => LD);
    
    v413: FDE1
        port map(Q0 => QI(7),
                 D0 => v139,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v414: FDE1
        port map(Q0 => QI(6),
                 D0 => v146,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v415: FDE1
        port map(Q0 => QI(5),
                 D0 => v142,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v416: AND2
        port map(Z0 => v130,
                 A0 => D6,
                 A1 => LD);
    
    v417: LXOR2
        port map(Z0 => v139,
                 A0 => v138,
                 A1 => v144);
    
    v418: AND2
        port map(Z0 => v140,
                 A0 => D7,
                 A1 => LD);
    
    v419: LXOR2
        port map(Z0 => v146,
                 A0 => v150,
                 A1 => v145);
    
    v420: LXOR2
        port map(Z0 => v142,
                 A0 => v141,
                 A1 => v148);
    
    v421: AND9
        port map(Z0 => v147,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v143,
                 A7 => CAI,
                 A8 => EN);
    
    v422: INV
        port map(ZN0 => v159,
                 A0 => LD);
    
    v423: AND2
        port map(Z0 => v157,
                 A0 => QI(9),
                 A1 => v159);
    
    v424: OR2
        port map(Z0 => v164,
                 A0 => v153,
                 A1 => v165);
    
    v425: AND2
        port map(Z0 => v166,
                 A0 => QI(10),
                 A1 => v159);
    
    v426: OR2
        port map(Z0 => v161,
                 A0 => v151,
                 A1 => v163);
    
    v427: AND2
        port map(Z0 => v154,
                 A0 => QI(11),
                 A1 => v159);
    
    v428: OR2
        port map(Z0 => v160,
                 A0 => v156,
                 A1 => v152);
    
    v429: AND12
        port map(Z0 => v165,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v159,
                 A10 => CAI,
                 A11 => EN);
    
    v430: AND13
        port map(Z0 => v163,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v159,
                 A11 => CAI,
                 A12 => EN);
    
    v431: AND14
        port map(Z0 => v152,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v205(10),
                 A11 => v159,
                 A12 => CAI,
                 A13 => EN);
    
    v432: INV
        port map(ZN0 => v205(9),
                 A0 => QI(9));
    
    v433: INV
        port map(ZN0 => v205(10),
                 A0 => QI(10));
    
    v434: INV
        port map(ZN0 => v205(11),
                 A0 => QI(11));
    
    v435: AND2
        port map(Z0 => v153,
                 A0 => D9,
                 A1 => LD);
    
    v436: FDE1
        port map(Q0 => QI(11),
                 D0 => v155,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v437: FDE1
        port map(Q0 => QI(10),
                 D0 => v162,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v438: FDE1
        port map(Q0 => QI(9),
                 D0 => v158,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v439: AND2
        port map(Z0 => v151,
                 A0 => D10,
                 A1 => LD);
    
    v440: LXOR2
        port map(Z0 => v155,
                 A0 => v154,
                 A1 => v160);
    
    v441: AND2
        port map(Z0 => v156,
                 A0 => D11,
                 A1 => LD);
    
    v442: LXOR2
        port map(Z0 => v162,
                 A0 => v166,
                 A1 => v161);
    
    v443: LXOR2
        port map(Z0 => v158,
                 A0 => v157,
                 A1 => v164);
    
    v444: INV
        port map(ZN0 => v167,
                 A0 => LD);
    
    v445: AND2
        port map(Z0 => v172,
                 A0 => QI(12),
                 A1 => v167);
    
    v446: OR2
        port map(Z0 => v176,
                 A0 => v171,
                 A1 => v177);
    
    v447: AND2
        port map(Z0 => v169,
                 A0 => QI(13),
                 A1 => v167);
    
    v448: OR2
        port map(Z0 => v174,
                 A0 => v168,
                 A1 => v175);
    
    v449: AND15
        port map(Z0 => v177,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v205(10),
                 A11 => v205(11),
                 A12 => v167,
                 A13 => CAI,
                 A14 => EN);
    
    v450: AND16
        port map(Z0 => v175,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v205(10),
                 A11 => v205(11),
                 A12 => v205(12),
                 A13 => v167,
                 A14 => CAI,
                 A15 => EN);
    
    v451: INV
        port map(ZN0 => v205(12),
                 A0 => QI(12));
    
    v452: INV
        port map(ZN0 => v205(13),
                 A0 => QI(13));
    
    v453: AND2
        port map(Z0 => v168,
                 A0 => D13,
                 A1 => LD);
    
    v454: AND2
        port map(Z0 => v171,
                 A0 => D12,
                 A1 => LD);
    
    v455: FDE1
        port map(Q0 => QI(13),
                 D0 => v170,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v456: FDE1
        port map(Q0 => QI(12),
                 D0 => v173,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v457: LXOR2
        port map(Z0 => v170,
                 A0 => v169,
                 A1 => v174);
    
    v458: LXOR2
        port map(Z0 => v173,
                 A0 => v172,
                 A1 => v176);
    
    v459: INV
        port map(ZN0 => v183,
                 A0 => LD);
    
    v460: AND2
        port map(Z0 => v188,
                 A0 => QI(14),
                 A1 => v183);
    
    v461: OR2
        port map(Z0 => v185,
                 A0 => v178,
                 A1 => v187);
    
    v462: AND2
        port map(Z0 => v180,
                 A0 => QI(15),
                 A1 => v183);
    
    v463: OR2
        port map(Z0 => v184,
                 A0 => v182,
                 A1 => v179);
    
    v464: AND17
        port map(Z0 => v187,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v205(10),
                 A11 => v205(11),
                 A12 => v205(12),
                 A13 => v205(13),
                 A14 => v183,
                 A15 => CAI,
                 A16 => EN);
    
    v465: AND18
        port map(Z0 => v179,
                 A0 => v205(0),
                 A1 => v205(1),
                 A2 => v205(2),
                 A3 => v205(3),
                 A4 => v205(4),
                 A5 => v205(5),
                 A6 => v205(6),
                 A7 => v205(7),
                 A8 => v205(8),
                 A9 => v205(9),
                 A10 => v205(10),
                 A11 => v205(11),
                 A12 => v205(12),
                 A13 => v205(13),
                 A14 => v205(14),
                 A15 => v183,
                 A16 => CAI,
                 A17 => EN);
    
    v466: INV
        port map(ZN0 => v205(14),
                 A0 => QI(14));
    
    v467: INV
        port map(ZN0 => v205(15),
                 A0 => QI(15));
    
    v468: FDE1
        port map(Q0 => QI(15),
                 D0 => v181,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v469: FDE1
        port map(Q0 => QI(14),
                 D0 => v186,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v470: AND2
        port map(Z0 => v178,
                 A0 => D14,
                 A1 => LD);
    
    v471: LXOR2
        port map(Z0 => v181,
                 A0 => v180,
                 A1 => v184);
    
    v472: AND2
        port map(Z0 => v182,
                 A0 => D15,
                 A1 => LD);
    
    v473: LXOR2
        port map(Z0 => v186,
                 A0 => v188,
                 A1 => v185);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBDA4 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBDA4;

architecture LATTICE_ARCH of CBDA4 is
    signal QI: std_logic_vector(0 to 3);
    signal v125: std_logic_vector(0 to 3);
    signal v116: std_logic;
    signal v104: std_logic;
    signal v102: std_logic;
    signal v112: std_logic;
    signal v111: std_logic;
    signal v103: std_logic;
    signal v113: std_logic;
    signal v120: std_logic;
    signal v118: std_logic;
    signal v105: std_logic;
    signal v117: std_logic;
    signal v115: std_logic;
    signal v114: std_logic;
    signal v110: std_logic;
    signal v107: std_logic;
    signal v119: std_logic;
    signal v106: std_logic;
    signal v108: std_logic;
    signal v109: std_logic;
    signal v100: std_logic;
    signal v101: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v160: FDE1
        port map(Q0 => QI(0),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v161: FDE1
        port map(Q0 => QI(1),
                 D0 => v118,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v162: AND2
        port map(Z0 => v100,
                 A0 => QI(0),
                 A1 => v116);
    
    v163: AND2
        port map(Z0 => v102,
                 A0 => D0,
                 A1 => LD);
    
    v164: AND2
        port map(Z0 => v105,
                 A0 => D1,
                 A1 => LD);
    
    v165: AND2
        port map(Z0 => v109,
                 A0 => QI(2),
                 A1 => v116);
    
    v166: AND2
        port map(Z0 => v108,
                 A0 => D2,
                 A1 => LD);
    
    v167: AND2
        port map(Z0 => v113,
                 A0 => QI(3),
                 A1 => v116);
    
    v168: AND2
        port map(Z0 => v112,
                 A0 => D3,
                 A1 => LD);
    
    v169: AND4
        port map(Z0 => v101,
                 A0 => v125(0),
                 A1 => CAI,
                 A2 => v116,
                 A3 => EN);
    
    v170: OR2
        port map(Z0 => v107,
                 A0 => v105,
                 A1 => v101);
    
    v171: OR2
        port map(Z0 => v110,
                 A0 => v108,
                 A1 => v111);
    
    v172: OR2
        port map(Z0 => v114,
                 A0 => v112,
                 A1 => v115);
    
    v173: AND5
        port map(Z0 => v111,
                 A0 => v125(0),
                 A1 => v125(1),
                 A2 => v116,
                 A3 => CAI,
                 A4 => EN);
    
    v174: AND6
        port map(Z0 => v115,
                 A0 => v125(0),
                 A1 => v125(1),
                 A2 => v125(2),
                 A3 => v116,
                 A4 => CAI,
                 A5 => EN);
    
    v175: AND2
        port map(Z0 => v106,
                 A0 => QI(1),
                 A1 => v116);
    
    v176: AND6
        port map(Z0 => CAO,
                 A0 => v125(0),
                 A1 => v125(1),
                 A2 => v125(2),
                 A3 => v125(3),
                 A4 => CAI,
                 A5 => EN);
    
    v177: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v178: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v179: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v180: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v181: AND3
        port map(Z0 => v103,
                 A0 => v116,
                 A1 => CAI,
                 A2 => EN);
    
    v182: INV
        port map(ZN0 => v125(0),
                 A0 => QI(0));
    
    v183: INV
        port map(ZN0 => v125(1),
                 A0 => QI(1));
    
    v184: INV
        port map(ZN0 => v125(2),
                 A0 => QI(2));
    
    v185: INV
        port map(ZN0 => v125(3),
                 A0 => QI(3));
    
    v186: FDE1
        port map(Q0 => QI(2),
                 D0 => v119,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v187: FDE1
        port map(Q0 => QI(3),
                 D0 => v120,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v188: LXOR2
        port map(Z0 => v117,
                 A0 => v100,
                 A1 => v104);
    
    v189: OR2
        port map(Z0 => v104,
                 A0 => v102,
                 A1 => v103);
    
    v190: LXOR2
        port map(Z0 => v118,
                 A0 => v106,
                 A1 => v107);
    
    v191: INV
        port map(ZN0 => v116,
                 A0 => LD);
    
    v192: LXOR2
        port map(Z0 => v119,
                 A0 => v109,
                 A1 => v110);
    
    v193: LXOR2
        port map(Z0 => v120,
                 A0 => v113,
                 A1 => v114);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBDA8 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBDA8;

architecture LATTICE_ARCH of CBDA8 is
    signal QI: std_logic_vector(0 to 7);
    signal v152: std_logic_vector(0 to 7);
    signal v118: std_logic;
    signal v106: std_logic;
    signal v124: std_logic;
    signal v104: std_logic;
    signal v114: std_logic;
    signal v133: std_logic;
    signal v113: std_logic;
    signal v105: std_logic;
    signal v115: std_logic;
    signal v122: std_logic;
    signal v120: std_logic;
    signal v107: std_logic;
    signal v137: std_logic;
    signal v119: std_logic;
    signal v117: std_logic;
    signal v143: std_logic;
    signal v116: std_logic;
    signal v112: std_logic;
    signal v109: std_logic;
    signal v121: std_logic;
    signal v108: std_logic;
    signal v110: std_logic;
    signal v111: std_logic;
    signal v102: std_logic;
    signal v123: std_logic;
    signal v127: std_logic;
    signal v134: std_logic;
    signal v128: std_logic;
    signal v103: std_logic;
    signal v138: std_logic;
    signal v129: std_logic;
    signal v139: std_logic;
    signal v130: std_logic;
    signal v135: std_logic;
    signal v125: std_logic;
    signal v140: std_logic;
    signal v131: std_logic;
    signal v126: std_logic;
    signal v132: std_logic;
    signal v141: std_logic;
    signal v136: std_logic;
    signal v142: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
begin
    v220: FDE1
        port map(Q0 => QI(0),
                 D0 => v119,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v221: FDE1
        port map(Q0 => QI(1),
                 D0 => v120,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v222: AND2
        port map(Z0 => v104,
                 A0 => D0,
                 A1 => LD);
    
    v223: AND3
        port map(Z0 => v105,
                 A0 => v118,
                 A1 => CAI,
                 A2 => EN);
    
    v224: AND2
        port map(Z0 => v107,
                 A0 => D1,
                 A1 => LD);
    
    v225: AND2
        port map(Z0 => v110,
                 A0 => D2,
                 A1 => LD);
    
    v226: AND2
        port map(Z0 => v114,
                 A0 => D3,
                 A1 => LD);
    
    v227: AND4
        port map(Z0 => v103,
                 A0 => v152(0),
                 A1 => CAI,
                 A2 => v118,
                 A3 => EN);
    
    v228: AND5
        port map(Z0 => v113,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v118,
                 A3 => CAI,
                 A4 => EN);
    
    v229: AND6
        port map(Z0 => v117,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v152(2),
                 A3 => v118,
                 A4 => CAI,
                 A5 => EN);
    
    v230: AND10
        port map(Z0 => CAO,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v152(2),
                 A3 => v152(3),
                 A4 => v152(4),
                 A5 => v152(5),
                 A6 => v152(6),
                 A7 => v152(7),
                 A8 => CAI,
                 A9 => EN);
    
    v231: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v232: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v233: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v234: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v235: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v236: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v237: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v238: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v239: OR2
        port map(Z0 => v106,
                 A0 => v104,
                 A1 => v105);
    
    v240: OR2
        port map(Z0 => v109,
                 A0 => v107,
                 A1 => v103);
    
    v241: OR2
        port map(Z0 => v112,
                 A0 => v110,
                 A1 => v113);
    
    v242: OR2
        port map(Z0 => v116,
                 A0 => v114,
                 A1 => v117);
    
    v243: AND2
        port map(Z0 => v102,
                 A0 => QI(0),
                 A1 => v118);
    
    v244: AND2
        port map(Z0 => v108,
                 A0 => QI(1),
                 A1 => v118);
    
    v245: AND2
        port map(Z0 => v111,
                 A0 => QI(2),
                 A1 => v118);
    
    v246: AND2
        port map(Z0 => v115,
                 A0 => QI(3),
                 A1 => v118);
    
    v247: INV
        port map(ZN0 => v152(0),
                 A0 => QI(0));
    
    v248: INV
        port map(ZN0 => v152(1),
                 A0 => QI(1));
    
    v249: INV
        port map(ZN0 => v152(2),
                 A0 => QI(2));
    
    v250: INV
        port map(ZN0 => v152(3),
                 A0 => QI(3));
    
    v251: FDE1
        port map(Q0 => QI(2),
                 D0 => v121,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v252: FDE1
        port map(Q0 => QI(3),
                 D0 => v122,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v253: LXOR2
        port map(Z0 => v119,
                 A0 => v102,
                 A1 => v106);
    
    v254: LXOR2
        port map(Z0 => v120,
                 A0 => v108,
                 A1 => v109);
    
    v255: INV
        port map(ZN0 => v118,
                 A0 => LD);
    
    v256: LXOR2
        port map(Z0 => v121,
                 A0 => v111,
                 A1 => v112);
    
    v257: LXOR2
        port map(Z0 => v122,
                 A0 => v115,
                 A1 => v116);
    
    v258: AND10
        port map(Z0 => v124,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v152(2),
                 A3 => v152(3),
                 A4 => v152(4),
                 A5 => v152(5),
                 A6 => v152(6),
                 A7 => v133,
                 A8 => CAI,
                 A9 => EN);
    
    v259: INV
        port map(ZN0 => v133,
                 A0 => LD);
    
    v260: OR2
        port map(Z0 => v141,
                 A0 => v131,
                 A1 => v142);
    
    v261: OR2
        port map(Z0 => v139,
                 A0 => v125,
                 A1 => v140);
    
    v262: OR2
        port map(Z0 => v136,
                 A0 => v123,
                 A1 => v138);
    
    v263: OR2
        port map(Z0 => v135,
                 A0 => v128,
                 A1 => v124);
    
    v264: AND2
        port map(Z0 => v132,
                 A0 => QI(4),
                 A1 => v133);
    
    v265: AND2
        port map(Z0 => v129,
                 A0 => QI(5),
                 A1 => v133);
    
    v266: AND2
        port map(Z0 => v143,
                 A0 => QI(6),
                 A1 => v133);
    
    v267: AND2
        port map(Z0 => v126,
                 A0 => QI(7),
                 A1 => v133);
    
    v268: INV
        port map(ZN0 => v152(4),
                 A0 => QI(4));
    
    v269: INV
        port map(ZN0 => v152(5),
                 A0 => QI(5));
    
    v270: INV
        port map(ZN0 => v152(6),
                 A0 => QI(6));
    
    v271: INV
        port map(ZN0 => v152(7),
                 A0 => QI(7));
    
    v272: AND7
        port map(Z0 => v142,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v152(2),
                 A3 => v152(3),
                 A4 => v133,
                 A5 => CAI,
                 A6 => EN);
    
    v273: AND8
        port map(Z0 => v140,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v152(2),
                 A3 => v152(3),
                 A4 => v152(4),
                 A5 => v133,
                 A6 => CAI,
                 A7 => EN);
    
    v274: AND2
        port map(Z0 => v125,
                 A0 => D5,
                 A1 => LD);
    
    v275: AND2
        port map(Z0 => v131,
                 A0 => D4,
                 A1 => LD);
    
    v276: FDE1
        port map(Q0 => QI(7),
                 D0 => v127,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v277: FDE1
        port map(Q0 => QI(6),
                 D0 => v137,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v278: FDE1
        port map(Q0 => QI(5),
                 D0 => v130,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v279: FDE1
        port map(Q0 => QI(4),
                 D0 => v134,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v280: AND2
        port map(Z0 => v123,
                 A0 => D6,
                 A1 => LD);
    
    v281: LXOR2
        port map(Z0 => v127,
                 A0 => v126,
                 A1 => v135);
    
    v282: AND2
        port map(Z0 => v128,
                 A0 => D7,
                 A1 => LD);
    
    v283: LXOR2
        port map(Z0 => v137,
                 A0 => v143,
                 A1 => v136);
    
    v284: LXOR2
        port map(Z0 => v130,
                 A0 => v129,
                 A1 => v139);
    
    v285: LXOR2
        port map(Z0 => v134,
                 A0 => v132,
                 A1 => v141);
    
    v286: AND9
        port map(Z0 => v138,
                 A0 => v152(0),
                 A1 => v152(1),
                 A2 => v152(2),
                 A3 => v152(3),
                 A4 => v152(4),
                 A5 => v152(5),
                 A6 => v133,
                 A7 => CAI,
                 A8 => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBDB4 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic;
         CS: IN std_logic);
end CBDB4;

architecture LATTICE_ARCH of CBDB4 is
    signal QI: std_logic_vector(0 to 3);
    signal v129: std_logic_vector(0 to 3);
    signal v119: std_logic;
    signal v107: std_logic;
    signal v105: std_logic;
    signal v115: std_logic;
    signal v120: std_logic;
    signal v106: std_logic;
    signal v116: std_logic;
    signal v124: std_logic;
    signal v122: std_logic;
    signal v108: std_logic;
    signal v121: std_logic;
    signal v118: std_logic;
    signal v109: std_logic;
    signal v117: std_logic;
    signal v114: std_logic;
    signal v111: std_logic;
    signal v123: std_logic;
    signal v110: std_logic;
    signal v112: std_logic;
    signal v113: std_logic;
    signal v103: std_logic;
    signal v104: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
begin
    v165: FDC1
        port map(Q0 => QI(0),
                 D0 => v121,
                 CLK => CLK,
                 SD => SD);
    
    v166: FDC1
        port map(Q0 => QI(1),
                 D0 => v122,
                 CLK => CLK,
                 SD => SD);
    
    v167: AND6
        port map(Z0 => v104,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => CAI,
                 A3 => v119,
                 A4 => EN,
                 A5 => v120);
    
    v168: AND7
        port map(Z0 => v118,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v119,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v120);
    
    v169: AND6
        port map(Z0 => CAO,
                 A0 => v129(0),
                 A1 => v129(1),
                 A2 => v129(2),
                 A3 => v129(3),
                 A4 => CAI,
                 A5 => EN);
    
    v170: INV
        port map(ZN0 => v120,
                 A0 => CS);
    
    v171: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v172: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v173: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v174: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v175: OR2
        port map(Z0 => v107,
                 A0 => v105,
                 A1 => v106);
    
    v176: OR2
        port map(Z0 => v111,
                 A0 => v108,
                 A1 => v109);
    
    v177: OR2
        port map(Z0 => v114,
                 A0 => v112,
                 A1 => v104);
    
    v178: OR2
        port map(Z0 => v117,
                 A0 => v115,
                 A1 => v118);
    
    v179: AND3
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => v119,
                 A2 => v120);
    
    v180: AND3
        port map(Z0 => v110,
                 A0 => QI(1),
                 A1 => v119,
                 A2 => v120);
    
    v181: AND3
        port map(Z0 => v113,
                 A0 => QI(2),
                 A1 => v119,
                 A2 => v120);
    
    v182: AND3
        port map(Z0 => v116,
                 A0 => QI(3),
                 A1 => v119,
                 A2 => v120);
    
    v183: INV
        port map(ZN0 => v129(0),
                 A0 => QI(0));
    
    v184: INV
        port map(ZN0 => v129(1),
                 A0 => QI(1));
    
    v185: INV
        port map(ZN0 => v129(2),
                 A0 => QI(2));
    
    v186: INV
        port map(ZN0 => v129(3),
                 A0 => QI(3));
    
    v187: FDC1
        port map(Q0 => QI(2),
                 D0 => v123,
                 CLK => CLK,
                 SD => SD);
    
    v188: FDC1
        port map(Q0 => QI(3),
                 D0 => v124,
                 CLK => CLK,
                 SD => SD);
    
    v189: AND3
        port map(Z0 => v105,
                 A0 => D0,
                 A1 => LD,
                 A2 => v120);
    
    v190: AND4
        port map(Z0 => v106,
                 A0 => v119,
                 A1 => CAI,
                 A2 => EN,
                 A3 => v120);
    
    v191: LXOR2
        port map(Z0 => v121,
                 A0 => v103,
                 A1 => v107);
    
    v192: LXOR2
        port map(Z0 => v122,
                 A0 => v110,
                 A1 => v111);
    
    v193: AND3
        port map(Z0 => v108,
                 A0 => D1,
                 A1 => LD,
                 A2 => v120);
    
    v194: INV
        port map(ZN0 => v119,
                 A0 => LD);
    
    v195: AND3
        port map(Z0 => v112,
                 A0 => D2,
                 A1 => LD,
                 A2 => v120);
    
    v196: LXOR2
        port map(Z0 => v123,
                 A0 => v113,
                 A1 => v114);
    
    v197: LXOR2
        port map(Z0 => v124,
                 A0 => v116,
                 A1 => v117);
    
    v198: AND3
        port map(Z0 => v115,
                 A0 => D3,
                 A1 => LD,
                 A2 => v120);
    
    v199: AND5
        port map(Z0 => v109,
                 A0 => v129(0),
                 A1 => CAI,
                 A2 => v119,
                 A3 => EN,
                 A4 => v120);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBDB8 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic;
         CS: IN std_logic);
end CBDB8;

architecture LATTICE_ARCH of CBDB8 is
    signal QI: std_logic_vector(0 to 7);
    signal v157: std_logic_vector(0 to 7);
    signal v121: std_logic;
    signal v109: std_logic;
    signal v128: std_logic;
    signal v107: std_logic;
    signal v117: std_logic;
    signal v130: std_logic;
    signal v122: std_logic;
    signal v108: std_logic;
    signal v141: std_logic;
    signal v118: std_logic;
    signal v139: std_logic;
    signal v126: std_logic;
    signal v124: std_logic;
    signal v110: std_logic;
    signal v147: std_logic;
    signal v140: std_logic;
    signal v123: std_logic;
    signal v120: std_logic;
    signal v111: std_logic;
    signal v131: std_logic;
    signal v119: std_logic;
    signal v116: std_logic;
    signal v113: std_logic;
    signal v134: std_logic;
    signal v132: std_logic;
    signal v125: std_logic;
    signal v112: std_logic;
    signal v145: std_logic;
    signal v136: std_logic;
    signal v138: std_logic;
    signal v114: std_logic;
    signal v148: std_logic;
    signal v142: std_logic;
    signal v129: std_logic;
    signal v143: std_logic;
    signal v135: std_logic;
    signal v115: std_logic;
    signal v146: std_logic;
    signal v137: std_logic;
    signal v144: std_logic;
    signal v133: std_logic;
    signal v105: std_logic;
    signal v106: std_logic;
    signal v127: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component AND11
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic);
    end component;
    for all : AND11 use entity LAT_VHD.AND11(LATTICE_ARCH);
    
begin
    v227: FDC1
        port map(Q0 => QI(0),
                 D0 => v123,
                 CLK => CLK,
                 SD => SD);
    
    v228: FDC1
        port map(Q0 => QI(1),
                 D0 => v124,
                 CLK => CLK,
                 SD => SD);
    
    v229: AND6
        port map(Z0 => v106,
                 A0 => v157(0),
                 A1 => v157(1),
                 A2 => CAI,
                 A3 => v121,
                 A4 => EN,
                 A5 => v122);
    
    v230: AND7
        port map(Z0 => v120,
                 A0 => v157(0),
                 A1 => v157(2),
                 A2 => v157(1),
                 A3 => v121,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v122);
    
    v231: AND10
        port map(Z0 => CAO,
                 A0 => v157(0),
                 A1 => v157(1),
                 A2 => v157(2),
                 A3 => v157(3),
                 A4 => v157(4),
                 A5 => v157(5),
                 A6 => v157(6),
                 A7 => v157(7),
                 A8 => CAI,
                 A9 => EN);
    
    v232: INV
        port map(ZN0 => v122,
                 A0 => CS);
    
    v233: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v234: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v235: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v236: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v237: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v238: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v239: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v240: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v241: OR2
        port map(Z0 => v119,
                 A0 => v117,
                 A1 => v120);
    
    v242: OR2
        port map(Z0 => v116,
                 A0 => v114,
                 A1 => v106);
    
    v243: OR2
        port map(Z0 => v113,
                 A0 => v110,
                 A1 => v111);
    
    v244: OR2
        port map(Z0 => v109,
                 A0 => v107,
                 A1 => v108);
    
    v245: AND3
        port map(Z0 => v105,
                 A0 => QI(0),
                 A1 => v121,
                 A2 => v122);
    
    v246: AND3
        port map(Z0 => v112,
                 A0 => QI(1),
                 A1 => v121,
                 A2 => v122);
    
    v247: AND3
        port map(Z0 => v115,
                 A0 => QI(2),
                 A1 => v121,
                 A2 => v122);
    
    v248: AND3
        port map(Z0 => v118,
                 A0 => QI(3),
                 A1 => v121,
                 A2 => v122);
    
    v249: INV
        port map(ZN0 => v157(0),
                 A0 => QI(0));
    
    v250: INV
        port map(ZN0 => v157(1),
                 A0 => QI(1));
    
    v251: INV
        port map(ZN0 => v157(2),
                 A0 => QI(2));
    
    v252: INV
        port map(ZN0 => v157(3),
                 A0 => QI(3));
    
    v253: FDC1
        port map(Q0 => QI(2),
                 D0 => v125,
                 CLK => CLK,
                 SD => SD);
    
    v254: FDC1
        port map(Q0 => QI(3),
                 D0 => v126,
                 CLK => CLK,
                 SD => SD);
    
    v255: AND3
        port map(Z0 => v107,
                 A0 => D0,
                 A1 => LD,
                 A2 => v122);
    
    v256: AND4
        port map(Z0 => v108,
                 A0 => v121,
                 A1 => CAI,
                 A2 => EN,
                 A3 => v122);
    
    v257: LXOR2
        port map(Z0 => v123,
                 A0 => v105,
                 A1 => v109);
    
    v258: LXOR2
        port map(Z0 => v124,
                 A0 => v112,
                 A1 => v113);
    
    v259: AND3
        port map(Z0 => v110,
                 A0 => D1,
                 A1 => LD,
                 A2 => v122);
    
    v260: INV
        port map(ZN0 => v121,
                 A0 => LD);
    
    v261: AND3
        port map(Z0 => v114,
                 A0 => D2,
                 A1 => LD,
                 A2 => v122);
    
    v262: LXOR2
        port map(Z0 => v125,
                 A0 => v115,
                 A1 => v116);
    
    v263: LXOR2
        port map(Z0 => v126,
                 A0 => v118,
                 A1 => v119);
    
    v264: AND3
        port map(Z0 => v117,
                 A0 => D3,
                 A1 => LD,
                 A2 => v122);
    
    v265: AND5
        port map(Z0 => v111,
                 A0 => v157(0),
                 A1 => CAI,
                 A2 => v121,
                 A3 => EN,
                 A4 => v122);
    
    v266: AND8
        port map(Z0 => v132,
                 A0 => v157(0),
                 A1 => v157(1),
                 A2 => v157(2),
                 A3 => v157(3),
                 A4 => v128,
                 A5 => CAI,
                 A6 => EN,
                 A7 => v141);
    
    v267: AND9
        port map(Z0 => v136,
                 A0 => v157(0),
                 A1 => v157(1),
                 A2 => v157(2),
                 A3 => v157(3),
                 A4 => v157(4),
                 A5 => v128,
                 A6 => CAI,
                 A7 => EN,
                 A8 => v141);
    
    v268: AND10
        port map(Z0 => v137,
                 A0 => v157(0),
                 A1 => v157(1),
                 A2 => v157(2),
                 A3 => v157(3),
                 A4 => v157(4),
                 A5 => v157(5),
                 A6 => v128,
                 A7 => CAI,
                 A8 => EN,
                 A9 => v141);
    
    v269: AND11
        port map(Z0 => v127,
                 A0 => v157(0),
                 A1 => v157(1),
                 A2 => v157(2),
                 A3 => v157(3),
                 A4 => v157(4),
                 A5 => v157(5),
                 A6 => v157(6),
                 A7 => v128,
                 A8 => CAI,
                 A9 => EN,
                 A10 => v141);
    
    v270: INV
        port map(ZN0 => v141,
                 A0 => CS);
    
    v271: OR2
        port map(Z0 => v129,
                 A0 => v131,
                 A1 => v132);
    
    v272: OR2
        port map(Z0 => v133,
                 A0 => v135,
                 A1 => v136);
    
    v273: OR2
        port map(Z0 => v140,
                 A0 => v138,
                 A1 => v137);
    
    v274: OR2
        port map(Z0 => v142,
                 A0 => v144,
                 A1 => v127);
    
    v275: AND3
        port map(Z0 => v130,
                 A0 => QI(4),
                 A1 => v128,
                 A2 => v141);
    
    v276: AND3
        port map(Z0 => v134,
                 A0 => QI(5),
                 A1 => v128,
                 A2 => v141);
    
    v277: AND3
        port map(Z0 => v139,
                 A0 => QI(6),
                 A1 => v128,
                 A2 => v141);
    
    v278: AND3
        port map(Z0 => v143,
                 A0 => QI(7),
                 A1 => v128,
                 A2 => v141);
    
    v279: INV
        port map(ZN0 => v157(4),
                 A0 => QI(4));
    
    v280: INV
        port map(ZN0 => v157(5),
                 A0 => QI(5));
    
    v281: INV
        port map(ZN0 => v157(6),
                 A0 => QI(6));
    
    v282: INV
        port map(ZN0 => v157(7),
                 A0 => QI(7));
    
    v283: INV
        port map(ZN0 => v128,
                 A0 => LD);
    
    v284: LXOR2
        port map(Z0 => v145,
                 A0 => v130,
                 A1 => v129);
    
    v285: FDC1
        port map(Q0 => QI(4),
                 D0 => v145,
                 CLK => CLK,
                 SD => SD);
    
    v286: AND3
        port map(Z0 => v131,
                 A0 => D4,
                 A1 => LD,
                 A2 => v141);
    
    v287: LXOR2
        port map(Z0 => v146,
                 A0 => v134,
                 A1 => v133);
    
    v288: FDC1
        port map(Q0 => QI(5),
                 D0 => v146,
                 CLK => CLK,
                 SD => SD);
    
    v289: AND3
        port map(Z0 => v135,
                 A0 => D5,
                 A1 => LD,
                 A2 => v141);
    
    v290: AND3
        port map(Z0 => v138,
                 A0 => D6,
                 A1 => LD,
                 A2 => v141);
    
    v291: FDC1
        port map(Q0 => QI(6),
                 D0 => v147,
                 CLK => CLK,
                 SD => SD);
    
    v292: LXOR2
        port map(Z0 => v147,
                 A0 => v139,
                 A1 => v140);
    
    v293: LXOR2
        port map(Z0 => v148,
                 A0 => v143,
                 A1 => v142);
    
    v294: FDC1
        port map(Q0 => QI(7),
                 D0 => v148,
                 CLK => CLK,
                 SD => SD);
    
    v295: AND3
        port map(Z0 => v144,
                 A0 => D7,
                 A1 => LD,
                 A2 => v141);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBU84 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic);
end CBU84;

architecture LATTICE_ARCH of CBU84 is
    signal QI: std_logic_vector(0 to 3);
    signal v103: std_logic;
    signal v110: std_logic;
    signal v108: std_logic;
    signal v107: std_logic;
    signal v106: std_logic;
    signal v105: std_logic;
    signal v104: std_logic;
    signal v109: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v128: FDC1
        port map(Q0 => QI(0),
                 D0 => v107,
                 CLK => CLK,
                 SD => SD);
    
    v129: FDC1
        port map(Q0 => QI(1),
                 D0 => v108,
                 CLK => CLK,
                 SD => SD);
    
    v130: AND2
        port map(Z0 => v103,
                 A0 => CAI,
                 A1 => EN);
    
    v131: AND3
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => EN);
    
    v132: AND4
        port map(Z0 => v105,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => CAI,
                 A3 => EN);
    
    v133: AND5
        port map(Z0 => v106,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => CAI,
                 A4 => EN);
    
    v134: AND6
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN);
    
    v135: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v136: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v137: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v138: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v139: FDC1
        port map(Q0 => QI(2),
                 D0 => v109,
                 CLK => CLK,
                 SD => SD);
    
    v140: FDC1
        port map(Q0 => QI(3),
                 D0 => v110,
                 CLK => CLK,
                 SD => SD);
    
    v141: LXOR2
        port map(Z0 => v107,
                 A0 => QI(0),
                 A1 => v103);
    
    v142: LXOR2
        port map(Z0 => v108,
                 A0 => QI(1),
                 A1 => v104);
    
    v143: LXOR2
        port map(Z0 => v109,
                 A0 => QI(2),
                 A1 => v105);
    
    v144: LXOR2
        port map(Z0 => v110,
                 A0 => QI(3),
                 A1 => v106);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBU88 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic);
end CBU88;

architecture LATTICE_ARCH of CBU88 is
    signal QI: std_logic_vector(0 to 7);
    signal v105: std_logic;
    signal v119: std_logic;
    signal v116: std_logic;
    signal v114: std_logic;
    signal v111: std_logic;
    signal v113: std_logic;
    signal v108: std_logic;
    signal v107: std_logic;
    signal v106: std_logic;
    signal v117: std_logic;
    signal v115: std_logic;
    signal v120: std_logic;
    signal v112: std_logic;
    signal v109: std_logic;
    signal v118: std_logic;
    signal v110: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v154: FDC1
        port map(Q0 => QI(0),
                 D0 => v113,
                 CLK => CLK,
                 SD => SD);
    
    v155: FDC1
        port map(Q0 => QI(1),
                 D0 => v114,
                 CLK => CLK,
                 SD => SD);
    
    v156: AND10
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => CAI,
                 A9 => EN);
    
    v157: AND2
        port map(Z0 => v105,
                 A0 => CAI,
                 A1 => EN);
    
    v158: AND3
        port map(Z0 => v106,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => EN);
    
    v159: AND4
        port map(Z0 => v107,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => CAI,
                 A3 => EN);
    
    v160: AND5
        port map(Z0 => v108,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => CAI,
                 A4 => EN);
    
    v161: AND6
        port map(Z0 => v109,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN);
    
    v162: AND7
        port map(Z0 => v110,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => CAI,
                 A6 => EN);
    
    v163: AND8
        port map(Z0 => v111,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => CAI,
                 A7 => EN);
    
    v164: AND9
        port map(Z0 => v112,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => CAI,
                 A8 => EN);
    
    v165: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v166: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v167: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v168: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v169: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v170: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v171: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v172: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v173: FDC1
        port map(Q0 => QI(2),
                 D0 => v115,
                 CLK => CLK,
                 SD => SD);
    
    v174: FDC1
        port map(Q0 => QI(3),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD);
    
    v175: LXOR2
        port map(Z0 => v113,
                 A0 => QI(0),
                 A1 => v105);
    
    v176: LXOR2
        port map(Z0 => v114,
                 A0 => QI(1),
                 A1 => v106);
    
    v177: LXOR2
        port map(Z0 => v115,
                 A0 => QI(2),
                 A1 => v107);
    
    v178: LXOR2
        port map(Z0 => v116,
                 A0 => QI(3),
                 A1 => v108);
    
    v179: LXOR2
        port map(Z0 => v117,
                 A0 => QI(4),
                 A1 => v109);
    
    v180: FDC1
        port map(Q0 => QI(4),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD);
    
    v181: LXOR2
        port map(Z0 => v118,
                 A0 => QI(5),
                 A1 => v110);
    
    v182: FDC1
        port map(Q0 => QI(5),
                 D0 => v118,
                 CLK => CLK,
                 SD => SD);
    
    v183: FDC1
        port map(Q0 => QI(6),
                 D0 => v119,
                 CLK => CLK,
                 SD => SD);
    
    v184: LXOR2
        port map(Z0 => v119,
                 A0 => QI(6),
                 A1 => v111);
    
    v185: LXOR2
        port map(Z0 => v120,
                 A0 => QI(7),
                 A1 => v112);
    
    v186: FDC1
        port map(Q0 => QI(7),
                 D0 => v120,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBU94 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBU94;

architecture LATTICE_ARCH of CBU94 is
    signal QI: std_logic_vector(0 to 3);
    signal v100: std_logic;
    signal v107: std_logic;
    signal v105: std_logic;
    signal v104: std_logic;
    signal v103: std_logic;
    signal v102: std_logic;
    signal v101: std_logic;
    signal v106: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v125: FDE1
        port map(Q0 => QI(0),
                 D0 => v104,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v126: FDE1
        port map(Q0 => QI(1),
                 D0 => v105,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v127: AND2
        port map(Z0 => v100,
                 A0 => CAI,
                 A1 => EN);
    
    v128: AND3
        port map(Z0 => v101,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => EN);
    
    v129: AND4
        port map(Z0 => v102,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => CAI,
                 A3 => EN);
    
    v130: AND5
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => CAI,
                 A4 => EN);
    
    v131: AND6
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN);
    
    v132: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v133: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v134: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v135: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v136: FDE1
        port map(Q0 => QI(2),
                 D0 => v106,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v137: FDE1
        port map(Q0 => QI(3),
                 D0 => v107,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v138: LXOR2
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => v100);
    
    v139: LXOR2
        port map(Z0 => v105,
                 A0 => QI(1),
                 A1 => v101);
    
    v140: LXOR2
        port map(Z0 => v106,
                 A0 => QI(2),
                 A1 => v102);
    
    v141: LXOR2
        port map(Z0 => v107,
                 A0 => QI(3),
                 A1 => v103);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBU98 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBU98;

architecture LATTICE_ARCH of CBU98 is
    signal QI: std_logic_vector(0 to 7);
    signal v102: std_logic;
    signal v116: std_logic;
    signal v113: std_logic;
    signal v111: std_logic;
    signal v108: std_logic;
    signal v110: std_logic;
    signal v105: std_logic;
    signal v104: std_logic;
    signal v103: std_logic;
    signal v114: std_logic;
    signal v112: std_logic;
    signal v117: std_logic;
    signal v109: std_logic;
    signal v106: std_logic;
    signal v115: std_logic;
    signal v107: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
begin
    v151: FDE1
        port map(Q0 => QI(0),
                 D0 => v110,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v152: FDE1
        port map(Q0 => QI(1),
                 D0 => v111,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v153: AND10
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => CAI,
                 A9 => EN);
    
    v154: AND2
        port map(Z0 => v102,
                 A0 => CAI,
                 A1 => EN);
    
    v155: AND3
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => EN);
    
    v156: AND4
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => CAI,
                 A3 => EN);
    
    v157: AND5
        port map(Z0 => v105,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => CAI,
                 A4 => EN);
    
    v158: AND6
        port map(Z0 => v106,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN);
    
    v159: AND7
        port map(Z0 => v107,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => CAI,
                 A6 => EN);
    
    v160: AND8
        port map(Z0 => v108,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => CAI,
                 A7 => EN);
    
    v161: AND9
        port map(Z0 => v109,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => CAI,
                 A8 => EN);
    
    v162: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v163: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v164: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v165: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v166: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v167: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v168: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v169: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v170: FDE1
        port map(Q0 => QI(2),
                 D0 => v112,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v171: FDE1
        port map(Q0 => QI(3),
                 D0 => v113,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v172: LXOR2
        port map(Z0 => v110,
                 A0 => QI(0),
                 A1 => v102);
    
    v173: LXOR2
        port map(Z0 => v111,
                 A0 => QI(1),
                 A1 => v103);
    
    v174: LXOR2
        port map(Z0 => v112,
                 A0 => QI(2),
                 A1 => v104);
    
    v175: LXOR2
        port map(Z0 => v113,
                 A0 => QI(3),
                 A1 => v105);
    
    v176: LXOR2
        port map(Z0 => v114,
                 A0 => QI(4),
                 A1 => v106);
    
    v177: FDE1
        port map(Q0 => QI(4),
                 D0 => v114,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v178: LXOR2
        port map(Z0 => v115,
                 A0 => QI(5),
                 A1 => v107);
    
    v179: FDE1
        port map(Q0 => QI(5),
                 D0 => v115,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v180: FDE1
        port map(Q0 => QI(6),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v181: LXOR2
        port map(Z0 => v116,
                 A0 => QI(6),
                 A1 => v108);
    
    v182: LXOR2
        port map(Z0 => v117,
                 A0 => QI(7),
                 A1 => v109);
    
    v183: FDE1
        port map(Q0 => QI(7),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUA16 is
    port(CAI: IN std_logic;
         CAO: OUT std_logic;
         CD: IN std_logic;
         CLK: IN std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D10: IN std_logic;
         D11: IN std_logic;
         D12: IN std_logic;
         D13: IN std_logic;
         D14: IN std_logic;
         D15: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         D8: IN std_logic;
         D9: IN std_logic;
         EN: IN std_logic;
         LD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q10: OUT std_logic;
         Q11: OUT std_logic;
         Q12: OUT std_logic;
         Q13: OUT std_logic;
         Q14: OUT std_logic;
         Q15: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         Q8: OUT std_logic;
         Q9: OUT std_logic;
         SD: IN std_logic);
end CBUA16;

architecture LATTICE_ARCH of CBUA16 is
    signal QI: std_logic_vector(0 to 15);
    signal v125: std_logic;
    signal v113: std_logic;
    signal v136: std_logic;
    signal v111: std_logic;
    signal v152: std_logic;
    signal v133: std_logic;
    signal v121: std_logic;
    signal v143: std_logic;
    signal v135: std_logic;
    signal v120: std_logic;
    signal v112: std_logic;
    signal v179: std_logic;
    signal v159: std_logic;
    signal v122: std_logic;
    signal v129: std_logic;
    signal v127: std_logic;
    signal v114: std_logic;
    signal v183: std_logic;
    signal v146: std_logic;
    signal v126: std_logic;
    signal v124: std_logic;
    signal v162: std_logic;
    signal v150: std_logic;
    signal v134: std_logic;
    signal v123: std_logic;
    signal v119: std_logic;
    signal v116: std_logic;
    signal v166: std_logic;
    signal v131: std_logic;
    signal v128: std_logic;
    signal v115: std_logic;
    signal v186: std_logic;
    signal v167: std_logic;
    signal v132: std_logic;
    signal v188: std_logic;
    signal v117: std_logic;
    signal v118: std_logic;
    signal v110: std_logic;
    signal v104: std_logic;
    signal v130: std_logic;
    signal v151: std_logic;
    signal v139: std_logic;
    signal v178: std_logic;
    signal v155: std_logic;
    signal v140: std_logic;
    signal v156: std_logic;
    signal v181: std_logic;
    signal v173: std_logic;
    signal v105: std_logic;
    signal v182: std_logic;
    signal v147: std_logic;
    signal v106: std_logic;
    signal v163: std_logic;
    signal v141: std_logic;
    signal v107: std_logic;
    signal v157: std_logic;
    signal v148: std_logic;
    signal v142: std_logic;
    signal v108: std_logic;
    signal v187: std_logic;
    signal v169: std_logic;
    signal v164: std_logic;
    signal v158: std_logic;
    signal v144: std_logic;
    signal v137: std_logic;
    signal v174: std_logic;
    signal v170: std_logic;
    signal v160: std_logic;
    signal v153: std_logic;
    signal v149: std_logic;
    signal v138: std_logic;
    signal v109: std_logic;
    signal v168: std_logic;
    signal v165: std_logic;
    signal v154: std_logic;
    signal v184: std_logic;
    signal v175: std_logic;
    signal v171: std_logic;
    signal v180: std_logic;
    signal v172: std_logic;
    signal v145: std_logic;
    signal v176: std_logic;
    signal v161: std_logic;
    signal v185: std_logic;
    signal v177: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND18
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic;
             A15: IN std_logic;
             A16: IN std_logic;
             A17: IN std_logic);
    end component;
    for all : AND18 use entity LAT_VHD.AND18(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND11
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic);
    end component;
    for all : AND11 use entity LAT_VHD.AND11(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component AND12
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic);
    end component;
    for all : AND12 use entity LAT_VHD.AND12(LATTICE_ARCH);
    
    component AND13
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic);
    end component;
    for all : AND13 use entity LAT_VHD.AND13(LATTICE_ARCH);
    
    component AND14
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic);
    end component;
    for all : AND14 use entity LAT_VHD.AND14(LATTICE_ARCH);
    
    component AND15
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic);
    end component;
    for all : AND15 use entity LAT_VHD.AND15(LATTICE_ARCH);
    
    component AND16
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic;
             A15: IN std_logic);
    end component;
    for all : AND16 use entity LAT_VHD.AND16(LATTICE_ARCH);
    
    component AND17
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic;
             A12: IN std_logic;
             A13: IN std_logic;
             A14: IN std_logic;
             A15: IN std_logic;
             A16: IN std_logic);
    end component;
    for all : AND17 use entity LAT_VHD.AND17(LATTICE_ARCH);
    
begin
    v307: FDE1
        port map(Q0 => QI(0),
                 D0 => v126,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v308: FDE1
        port map(Q0 => QI(1),
                 D0 => v127,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v309: AND2
        port map(Z0 => v111,
                 A0 => D0,
                 A1 => LD);
    
    v310: AND3
        port map(Z0 => v112,
                 A0 => v125,
                 A1 => CAI,
                 A2 => EN);
    
    v311: AND2
        port map(Z0 => v114,
                 A0 => D1,
                 A1 => LD);
    
    v312: AND2
        port map(Z0 => v117,
                 A0 => D2,
                 A1 => LD);
    
    v313: AND2
        port map(Z0 => v121,
                 A0 => D3,
                 A1 => LD);
    
    v314: AND4
        port map(Z0 => v105,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v125,
                 A3 => EN);
    
    v315: AND5
        port map(Z0 => v120,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => v125,
                 A3 => CAI,
                 A4 => EN);
    
    v316: AND6
        port map(Z0 => v124,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v125,
                 A4 => CAI,
                 A5 => EN);
    
    v317: AND18
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => QI(10),
                 A11 => QI(11),
                 A12 => QI(12),
                 A13 => QI(13),
                 A14 => QI(14),
                 A15 => QI(15),
                 A16 => CAI,
                 A17 => EN);
    
    v318: AND2
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => v125);
    
    v319: OR2
        port map(Z0 => v113,
                 A0 => v111,
                 A1 => v112);
    
    v320: BUF
        port map(Z0 => Q15,
                 A0 => QI(15));
    
    v321: BUF
        port map(Z0 => Q11,
                 A0 => QI(11));
    
    v322: BUF
        port map(Z0 => Q9,
                 A0 => QI(9));
    
    v323: BUF
        port map(Z0 => Q8,
                 A0 => QI(8));
    
    v324: BUF
        port map(Z0 => Q14,
                 A0 => QI(14));
    
    v325: BUF
        port map(Z0 => Q13,
                 A0 => QI(13));
    
    v326: BUF
        port map(Z0 => Q12,
                 A0 => QI(12));
    
    v327: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v328: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v329: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v330: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v331: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v332: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v333: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v334: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v335: BUF
        port map(Z0 => Q10,
                 A0 => QI(10));
    
    v336: AND2
        port map(Z0 => v115,
                 A0 => QI(1),
                 A1 => v125);
    
    v337: OR2
        port map(Z0 => v116,
                 A0 => v114,
                 A1 => v105);
    
    v338: AND2
        port map(Z0 => v118,
                 A0 => QI(2),
                 A1 => v125);
    
    v339: OR2
        port map(Z0 => v119,
                 A0 => v117,
                 A1 => v120);
    
    v340: AND2
        port map(Z0 => v122,
                 A0 => QI(3),
                 A1 => v125);
    
    v341: OR2
        port map(Z0 => v123,
                 A0 => v121,
                 A1 => v124);
    
    v342: OR2
        port map(Z0 => v110,
                 A0 => v106,
                 A1 => v108);
    
    v343: AND2
        port map(Z0 => v109,
                 A0 => QI(4),
                 A1 => v125);
    
    v344: LXOR2
        port map(Z0 => v107,
                 A0 => v109,
                 A1 => v110);
    
    v345: FDE1
        port map(Q0 => QI(4),
                 D0 => v107,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v346: AND2
        port map(Z0 => v106,
                 A0 => D4,
                 A1 => LD);
    
    v347: AND7
        port map(Z0 => v108,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => v125,
                 A5 => CAI,
                 A6 => EN);
    
    v348: FDE1
        port map(Q0 => QI(2),
                 D0 => v128,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v349: FDE1
        port map(Q0 => QI(3),
                 D0 => v129,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v350: LXOR2
        port map(Z0 => v126,
                 A0 => v104,
                 A1 => v113);
    
    v351: LXOR2
        port map(Z0 => v127,
                 A0 => v115,
                 A1 => v116);
    
    v352: INV
        port map(ZN0 => v125,
                 A0 => LD);
    
    v353: LXOR2
        port map(Z0 => v128,
                 A0 => v118,
                 A1 => v119);
    
    v354: LXOR2
        port map(Z0 => v129,
                 A0 => v122,
                 A1 => v123);
    
    v355: AND10
        port map(Z0 => v136,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => v143,
                 A8 => CAI,
                 A9 => EN);
    
    v356: INV
        port map(ZN0 => v143,
                 A0 => LD);
    
    v357: AND2
        port map(Z0 => v141,
                 A0 => QI(5),
                 A1 => v143);
    
    v358: OR2
        port map(Z0 => v148,
                 A0 => v137,
                 A1 => v149);
    
    v359: AND2
        port map(Z0 => v150,
                 A0 => QI(6),
                 A1 => v143);
    
    v360: OR2
        port map(Z0 => v145,
                 A0 => v130,
                 A1 => v147);
    
    v361: AND2
        port map(Z0 => v138,
                 A0 => QI(7),
                 A1 => v143);
    
    v362: OR2
        port map(Z0 => v144,
                 A0 => v140,
                 A1 => v136);
    
    v363: OR2
        port map(Z0 => v134,
                 A0 => v131,
                 A1 => v135);
    
    v364: AND2
        port map(Z0 => v133,
                 A0 => QI(8),
                 A1 => v143);
    
    v365: LXOR2
        port map(Z0 => v132,
                 A0 => v133,
                 A1 => v134);
    
    v366: AND2
        port map(Z0 => v131,
                 A0 => D8,
                 A1 => LD);
    
    v367: FDE1
        port map(Q0 => QI(8),
                 D0 => v132,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v368: AND11
        port map(Z0 => v135,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => v143,
                 A9 => CAI,
                 A10 => EN);
    
    v369: AND8
        port map(Z0 => v149,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => v143,
                 A6 => CAI,
                 A7 => EN);
    
    v370: AND2
        port map(Z0 => v137,
                 A0 => D5,
                 A1 => LD);
    
    v371: FDE1
        port map(Q0 => QI(7),
                 D0 => v139,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v372: FDE1
        port map(Q0 => QI(6),
                 D0 => v146,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v373: FDE1
        port map(Q0 => QI(5),
                 D0 => v142,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v374: AND2
        port map(Z0 => v130,
                 A0 => D6,
                 A1 => LD);
    
    v375: LXOR2
        port map(Z0 => v139,
                 A0 => v138,
                 A1 => v144);
    
    v376: AND2
        port map(Z0 => v140,
                 A0 => D7,
                 A1 => LD);
    
    v377: LXOR2
        port map(Z0 => v146,
                 A0 => v150,
                 A1 => v145);
    
    v378: LXOR2
        port map(Z0 => v142,
                 A0 => v141,
                 A1 => v148);
    
    v379: AND9
        port map(Z0 => v147,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => v143,
                 A7 => CAI,
                 A8 => EN);
    
    v380: INV
        port map(ZN0 => v159,
                 A0 => LD);
    
    v381: AND2
        port map(Z0 => v157,
                 A0 => QI(9),
                 A1 => v159);
    
    v382: OR2
        port map(Z0 => v164,
                 A0 => v153,
                 A1 => v165);
    
    v383: AND2
        port map(Z0 => v166,
                 A0 => QI(10),
                 A1 => v159);
    
    v384: OR2
        port map(Z0 => v161,
                 A0 => v151,
                 A1 => v163);
    
    v385: AND2
        port map(Z0 => v154,
                 A0 => QI(11),
                 A1 => v159);
    
    v386: OR2
        port map(Z0 => v160,
                 A0 => v156,
                 A1 => v152);
    
    v387: AND12
        port map(Z0 => v165,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => v159,
                 A10 => CAI,
                 A11 => EN);
    
    v388: AND13
        port map(Z0 => v163,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => v159,
                 A11 => CAI,
                 A12 => EN);
    
    v389: AND14
        port map(Z0 => v152,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => QI(10),
                 A11 => v159,
                 A12 => CAI,
                 A13 => EN);
    
    v390: AND2
        port map(Z0 => v153,
                 A0 => D9,
                 A1 => LD);
    
    v391: FDE1
        port map(Q0 => QI(11),
                 D0 => v155,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v392: FDE1
        port map(Q0 => QI(10),
                 D0 => v162,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v393: FDE1
        port map(Q0 => QI(9),
                 D0 => v158,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v394: AND2
        port map(Z0 => v151,
                 A0 => D10,
                 A1 => LD);
    
    v395: LXOR2
        port map(Z0 => v155,
                 A0 => v154,
                 A1 => v160);
    
    v396: AND2
        port map(Z0 => v156,
                 A0 => D11,
                 A1 => LD);
    
    v397: LXOR2
        port map(Z0 => v162,
                 A0 => v166,
                 A1 => v161);
    
    v398: LXOR2
        port map(Z0 => v158,
                 A0 => v157,
                 A1 => v164);
    
    v399: INV
        port map(ZN0 => v167,
                 A0 => LD);
    
    v400: AND2
        port map(Z0 => v172,
                 A0 => QI(12),
                 A1 => v167);
    
    v401: OR2
        port map(Z0 => v176,
                 A0 => v171,
                 A1 => v177);
    
    v402: AND2
        port map(Z0 => v169,
                 A0 => QI(13),
                 A1 => v167);
    
    v403: OR2
        port map(Z0 => v174,
                 A0 => v168,
                 A1 => v175);
    
    v404: AND15
        port map(Z0 => v177,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => QI(10),
                 A11 => QI(11),
                 A12 => v167,
                 A13 => CAI,
                 A14 => EN);
    
    v405: AND16
        port map(Z0 => v175,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => QI(10),
                 A11 => QI(11),
                 A12 => QI(12),
                 A13 => v167,
                 A14 => CAI,
                 A15 => EN);
    
    v406: AND2
        port map(Z0 => v168,
                 A0 => D13,
                 A1 => LD);
    
    v407: AND2
        port map(Z0 => v171,
                 A0 => D12,
                 A1 => LD);
    
    v408: FDE1
        port map(Q0 => QI(13),
                 D0 => v170,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v409: FDE1
        port map(Q0 => QI(12),
                 D0 => v173,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v410: LXOR2
        port map(Z0 => v170,
                 A0 => v169,
                 A1 => v174);
    
    v411: LXOR2
        port map(Z0 => v173,
                 A0 => v172,
                 A1 => v176);
    
    v412: INV
        port map(ZN0 => v183,
                 A0 => LD);
    
    v413: AND2
        port map(Z0 => v188,
                 A0 => QI(14),
                 A1 => v183);
    
    v414: OR2
        port map(Z0 => v185,
                 A0 => v178,
                 A1 => v187);
    
    v415: AND2
        port map(Z0 => v180,
                 A0 => QI(15),
                 A1 => v183);
    
    v416: OR2
        port map(Z0 => v184,
                 A0 => v182,
                 A1 => v179);
    
    v417: AND17
        port map(Z0 => v187,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => QI(10),
                 A11 => QI(11),
                 A12 => QI(12),
                 A13 => QI(13),
                 A14 => v183,
                 A15 => CAI,
                 A16 => EN);
    
    v418: AND18
        port map(Z0 => v179,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => QI(8),
                 A9 => QI(9),
                 A10 => QI(10),
                 A11 => QI(11),
                 A12 => QI(12),
                 A13 => QI(13),
                 A14 => QI(14),
                 A15 => v183,
                 A16 => CAI,
                 A17 => EN);
    
    v419: FDE1
        port map(Q0 => QI(15),
                 D0 => v181,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v420: FDE1
        port map(Q0 => QI(14),
                 D0 => v186,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v421: AND2
        port map(Z0 => v178,
                 A0 => D14,
                 A1 => LD);
    
    v422: LXOR2
        port map(Z0 => v181,
                 A0 => v180,
                 A1 => v184);
    
    v423: AND2
        port map(Z0 => v182,
                 A0 => D15,
                 A1 => LD);
    
    v424: LXOR2
        port map(Z0 => v186,
                 A0 => v188,
                 A1 => v185);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUA4 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBUA4;

architecture LATTICE_ARCH of CBUA4 is
    signal QI: std_logic_vector(0 to 3);
    signal v116: std_logic;
    signal v104: std_logic;
    signal v102: std_logic;
    signal v112: std_logic;
    signal v111: std_logic;
    signal v103: std_logic;
    signal v113: std_logic;
    signal v120: std_logic;
    signal v118: std_logic;
    signal v105: std_logic;
    signal v117: std_logic;
    signal v115: std_logic;
    signal v114: std_logic;
    signal v110: std_logic;
    signal v107: std_logic;
    signal v119: std_logic;
    signal v106: std_logic;
    signal v108: std_logic;
    signal v109: std_logic;
    signal v100: std_logic;
    signal v101: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
begin
    v151: FDE1
        port map(Q0 => QI(0),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v152: FDE1
        port map(Q0 => QI(1),
                 D0 => v118,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v153: AND2
        port map(Z0 => v100,
                 A0 => QI(0),
                 A1 => v116);
    
    v154: AND2
        port map(Z0 => v102,
                 A0 => D0,
                 A1 => LD);
    
    v155: AND2
        port map(Z0 => v105,
                 A0 => D1,
                 A1 => LD);
    
    v156: AND2
        port map(Z0 => v109,
                 A0 => QI(2),
                 A1 => v116);
    
    v157: AND2
        port map(Z0 => v108,
                 A0 => D2,
                 A1 => LD);
    
    v158: AND2
        port map(Z0 => v113,
                 A0 => QI(3),
                 A1 => v116);
    
    v159: AND2
        port map(Z0 => v112,
                 A0 => D3,
                 A1 => LD);
    
    v160: AND4
        port map(Z0 => v101,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v116,
                 A3 => EN);
    
    v161: OR2
        port map(Z0 => v107,
                 A0 => v105,
                 A1 => v101);
    
    v162: OR2
        port map(Z0 => v110,
                 A0 => v108,
                 A1 => v111);
    
    v163: OR2
        port map(Z0 => v114,
                 A0 => v112,
                 A1 => v115);
    
    v164: AND5
        port map(Z0 => v111,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => v116,
                 A3 => CAI,
                 A4 => EN);
    
    v165: AND6
        port map(Z0 => v115,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v116,
                 A4 => CAI,
                 A5 => EN);
    
    v166: AND2
        port map(Z0 => v106,
                 A0 => QI(1),
                 A1 => v116);
    
    v167: AND6
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN);
    
    v168: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v169: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v170: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v171: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v172: AND3
        port map(Z0 => v103,
                 A0 => v116,
                 A1 => CAI,
                 A2 => EN);
    
    v173: FDE1
        port map(Q0 => QI(2),
                 D0 => v119,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v174: FDE1
        port map(Q0 => QI(3),
                 D0 => v120,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v175: LXOR2
        port map(Z0 => v117,
                 A0 => v100,
                 A1 => v104);
    
    v176: OR2
        port map(Z0 => v104,
                 A0 => v102,
                 A1 => v103);
    
    v177: LXOR2
        port map(Z0 => v118,
                 A0 => v106,
                 A1 => v107);
    
    v178: INV
        port map(ZN0 => v116,
                 A0 => LD);
    
    v179: LXOR2
        port map(Z0 => v119,
                 A0 => v109,
                 A1 => v110);
    
    v180: LXOR2
        port map(Z0 => v120,
                 A0 => v113,
                 A1 => v114);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUA8 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end CBUA8;

architecture LATTICE_ARCH of CBUA8 is
    signal QI: std_logic_vector(0 to 7);
    signal v118: std_logic;
    signal v106: std_logic;
    signal v124: std_logic;
    signal v104: std_logic;
    signal v114: std_logic;
    signal v133: std_logic;
    signal v113: std_logic;
    signal v105: std_logic;
    signal v115: std_logic;
    signal v122: std_logic;
    signal v120: std_logic;
    signal v107: std_logic;
    signal v137: std_logic;
    signal v119: std_logic;
    signal v117: std_logic;
    signal v143: std_logic;
    signal v116: std_logic;
    signal v112: std_logic;
    signal v109: std_logic;
    signal v121: std_logic;
    signal v108: std_logic;
    signal v110: std_logic;
    signal v111: std_logic;
    signal v102: std_logic;
    signal v123: std_logic;
    signal v127: std_logic;
    signal v134: std_logic;
    signal v128: std_logic;
    signal v103: std_logic;
    signal v138: std_logic;
    signal v129: std_logic;
    signal v139: std_logic;
    signal v130: std_logic;
    signal v135: std_logic;
    signal v125: std_logic;
    signal v140: std_logic;
    signal v131: std_logic;
    signal v126: std_logic;
    signal v132: std_logic;
    signal v141: std_logic;
    signal v136: std_logic;
    signal v142: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
begin
    v203: FDE1
        port map(Q0 => QI(0),
                 D0 => v119,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v204: FDE1
        port map(Q0 => QI(1),
                 D0 => v120,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v205: AND2
        port map(Z0 => v104,
                 A0 => D0,
                 A1 => LD);
    
    v206: AND3
        port map(Z0 => v105,
                 A0 => v118,
                 A1 => CAI,
                 A2 => EN);
    
    v207: AND2
        port map(Z0 => v107,
                 A0 => D1,
                 A1 => LD);
    
    v208: AND2
        port map(Z0 => v110,
                 A0 => D2,
                 A1 => LD);
    
    v209: AND2
        port map(Z0 => v114,
                 A0 => D3,
                 A1 => LD);
    
    v210: AND4
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v118,
                 A3 => EN);
    
    v211: AND5
        port map(Z0 => v113,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => v118,
                 A3 => CAI,
                 A4 => EN);
    
    v212: AND6
        port map(Z0 => v117,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v118,
                 A4 => CAI,
                 A5 => EN);
    
    v213: AND10
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => CAI,
                 A9 => EN);
    
    v214: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v215: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v216: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v217: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v218: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v219: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v220: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v221: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v222: OR2
        port map(Z0 => v106,
                 A0 => v104,
                 A1 => v105);
    
    v223: OR2
        port map(Z0 => v109,
                 A0 => v107,
                 A1 => v103);
    
    v224: OR2
        port map(Z0 => v112,
                 A0 => v110,
                 A1 => v113);
    
    v225: OR2
        port map(Z0 => v116,
                 A0 => v114,
                 A1 => v117);
    
    v226: AND2
        port map(Z0 => v102,
                 A0 => QI(0),
                 A1 => v118);
    
    v227: AND2
        port map(Z0 => v108,
                 A0 => QI(1),
                 A1 => v118);
    
    v228: AND2
        port map(Z0 => v111,
                 A0 => QI(2),
                 A1 => v118);
    
    v229: AND2
        port map(Z0 => v115,
                 A0 => QI(3),
                 A1 => v118);
    
    v230: FDE1
        port map(Q0 => QI(2),
                 D0 => v121,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v231: FDE1
        port map(Q0 => QI(3),
                 D0 => v122,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v232: LXOR2
        port map(Z0 => v119,
                 A0 => v102,
                 A1 => v106);
    
    v233: LXOR2
        port map(Z0 => v120,
                 A0 => v108,
                 A1 => v109);
    
    v234: INV
        port map(ZN0 => v118,
                 A0 => LD);
    
    v235: LXOR2
        port map(Z0 => v121,
                 A0 => v111,
                 A1 => v112);
    
    v236: LXOR2
        port map(Z0 => v122,
                 A0 => v115,
                 A1 => v116);
    
    v237: AND10
        port map(Z0 => v124,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => v133,
                 A8 => CAI,
                 A9 => EN);
    
    v238: INV
        port map(ZN0 => v133,
                 A0 => LD);
    
    v239: OR2
        port map(Z0 => v141,
                 A0 => v131,
                 A1 => v142);
    
    v240: OR2
        port map(Z0 => v139,
                 A0 => v125,
                 A1 => v140);
    
    v241: OR2
        port map(Z0 => v136,
                 A0 => v123,
                 A1 => v138);
    
    v242: OR2
        port map(Z0 => v135,
                 A0 => v128,
                 A1 => v124);
    
    v243: AND2
        port map(Z0 => v132,
                 A0 => QI(4),
                 A1 => v133);
    
    v244: AND2
        port map(Z0 => v129,
                 A0 => QI(5),
                 A1 => v133);
    
    v245: AND2
        port map(Z0 => v143,
                 A0 => QI(6),
                 A1 => v133);
    
    v246: AND2
        port map(Z0 => v126,
                 A0 => QI(7),
                 A1 => v133);
    
    v247: AND7
        port map(Z0 => v142,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => v133,
                 A5 => CAI,
                 A6 => EN);
    
    v248: AND8
        port map(Z0 => v140,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => v133,
                 A6 => CAI,
                 A7 => EN);
    
    v249: AND2
        port map(Z0 => v125,
                 A0 => D5,
                 A1 => LD);
    
    v250: AND2
        port map(Z0 => v131,
                 A0 => D4,
                 A1 => LD);
    
    v251: FDE1
        port map(Q0 => QI(7),
                 D0 => v127,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v252: FDE1
        port map(Q0 => QI(6),
                 D0 => v137,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v253: FDE1
        port map(Q0 => QI(5),
                 D0 => v130,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v254: FDE1
        port map(Q0 => QI(4),
                 D0 => v134,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v255: AND2
        port map(Z0 => v123,
                 A0 => D6,
                 A1 => LD);
    
    v256: LXOR2
        port map(Z0 => v127,
                 A0 => v126,
                 A1 => v135);
    
    v257: AND2
        port map(Z0 => v128,
                 A0 => D7,
                 A1 => LD);
    
    v258: LXOR2
        port map(Z0 => v137,
                 A0 => v143,
                 A1 => v136);
    
    v259: LXOR2
        port map(Z0 => v130,
                 A0 => v129,
                 A1 => v139);
    
    v260: LXOR2
        port map(Z0 => v134,
                 A0 => v132,
                 A1 => v141);
    
    v261: AND9
        port map(Z0 => v138,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => v133,
                 A7 => CAI,
                 A8 => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUB4 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic;
         CS: IN std_logic);
end CBUB4;

architecture LATTICE_ARCH of CBUB4 is
    signal QI: std_logic_vector(0 to 3);
    signal v119: std_logic;
    signal v107: std_logic;
    signal v105: std_logic;
    signal v115: std_logic;
    signal v120: std_logic;
    signal v106: std_logic;
    signal v116: std_logic;
    signal v124: std_logic;
    signal v122: std_logic;
    signal v108: std_logic;
    signal v121: std_logic;
    signal v118: std_logic;
    signal v109: std_logic;
    signal v117: std_logic;
    signal v114: std_logic;
    signal v111: std_logic;
    signal v123: std_logic;
    signal v110: std_logic;
    signal v112: std_logic;
    signal v113: std_logic;
    signal v103: std_logic;
    signal v104: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
begin
    v156: FDC1
        port map(Q0 => QI(0),
                 D0 => v121,
                 CLK => CLK,
                 SD => SD);
    
    v157: FDC1
        port map(Q0 => QI(1),
                 D0 => v122,
                 CLK => CLK,
                 SD => SD);
    
    v158: AND6
        port map(Z0 => v104,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => CAI,
                 A3 => v119,
                 A4 => EN,
                 A5 => v120);
    
    v159: AND7
        port map(Z0 => v118,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v119,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v120);
    
    v160: AND6
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN);
    
    v161: INV
        port map(ZN0 => v120,
                 A0 => CS);
    
    v162: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v163: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v164: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v165: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v166: OR2
        port map(Z0 => v107,
                 A0 => v105,
                 A1 => v106);
    
    v167: OR2
        port map(Z0 => v111,
                 A0 => v108,
                 A1 => v109);
    
    v168: OR2
        port map(Z0 => v114,
                 A0 => v112,
                 A1 => v104);
    
    v169: OR2
        port map(Z0 => v117,
                 A0 => v115,
                 A1 => v118);
    
    v170: AND3
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => v119,
                 A2 => v120);
    
    v171: AND3
        port map(Z0 => v110,
                 A0 => QI(1),
                 A1 => v119,
                 A2 => v120);
    
    v172: AND3
        port map(Z0 => v113,
                 A0 => QI(2),
                 A1 => v119,
                 A2 => v120);
    
    v173: AND3
        port map(Z0 => v116,
                 A0 => QI(3),
                 A1 => v119,
                 A2 => v120);
    
    v174: FDC1
        port map(Q0 => QI(2),
                 D0 => v123,
                 CLK => CLK,
                 SD => SD);
    
    v175: FDC1
        port map(Q0 => QI(3),
                 D0 => v124,
                 CLK => CLK,
                 SD => SD);
    
    v176: AND3
        port map(Z0 => v105,
                 A0 => D0,
                 A1 => LD,
                 A2 => v120);
    
    v177: AND4
        port map(Z0 => v106,
                 A0 => v119,
                 A1 => CAI,
                 A2 => EN,
                 A3 => v120);
    
    v178: LXOR2
        port map(Z0 => v121,
                 A0 => v103,
                 A1 => v107);
    
    v179: LXOR2
        port map(Z0 => v122,
                 A0 => v110,
                 A1 => v111);
    
    v180: AND3
        port map(Z0 => v108,
                 A0 => D1,
                 A1 => LD,
                 A2 => v120);
    
    v181: INV
        port map(ZN0 => v119,
                 A0 => LD);
    
    v182: AND3
        port map(Z0 => v112,
                 A0 => D2,
                 A1 => LD,
                 A2 => v120);
    
    v183: LXOR2
        port map(Z0 => v123,
                 A0 => v113,
                 A1 => v114);
    
    v184: LXOR2
        port map(Z0 => v124,
                 A0 => v116,
                 A1 => v117);
    
    v185: AND3
        port map(Z0 => v115,
                 A0 => D3,
                 A1 => LD,
                 A2 => v120);
    
    v186: AND5
        port map(Z0 => v109,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v119,
                 A3 => EN,
                 A4 => v120);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUB8 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic;
         CS: IN std_logic);
end CBUB8;

architecture LATTICE_ARCH of CBUB8 is
    signal QI: std_logic_vector(0 to 7);
    signal v121: std_logic;
    signal v109: std_logic;
    signal v128: std_logic;
    signal v107: std_logic;
    signal v117: std_logic;
    signal v130: std_logic;
    signal v122: std_logic;
    signal v108: std_logic;
    signal v141: std_logic;
    signal v118: std_logic;
    signal v139: std_logic;
    signal v126: std_logic;
    signal v124: std_logic;
    signal v110: std_logic;
    signal v147: std_logic;
    signal v140: std_logic;
    signal v123: std_logic;
    signal v120: std_logic;
    signal v111: std_logic;
    signal v131: std_logic;
    signal v119: std_logic;
    signal v116: std_logic;
    signal v113: std_logic;
    signal v134: std_logic;
    signal v132: std_logic;
    signal v125: std_logic;
    signal v112: std_logic;
    signal v145: std_logic;
    signal v136: std_logic;
    signal v138: std_logic;
    signal v114: std_logic;
    signal v148: std_logic;
    signal v142: std_logic;
    signal v129: std_logic;
    signal v143: std_logic;
    signal v135: std_logic;
    signal v115: std_logic;
    signal v146: std_logic;
    signal v137: std_logic;
    signal v144: std_logic;
    signal v133: std_logic;
    signal v105: std_logic;
    signal v106: std_logic;
    signal v127: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component AND11
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic);
    end component;
    for all : AND11 use entity LAT_VHD.AND11(LATTICE_ARCH);
    
begin
    v210: FDC1
        port map(Q0 => QI(0),
                 D0 => v123,
                 CLK => CLK,
                 SD => SD);
    
    v211: FDC1
        port map(Q0 => QI(1),
                 D0 => v124,
                 CLK => CLK,
                 SD => SD);
    
    v212: AND6
        port map(Z0 => v106,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => CAI,
                 A3 => v121,
                 A4 => EN,
                 A5 => v122);
    
    v213: AND7
        port map(Z0 => v120,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v121,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v122);
    
    v214: AND10
        port map(Z0 => CAO,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => CAI,
                 A9 => EN);
    
    v215: INV
        port map(ZN0 => v122,
                 A0 => CS);
    
    v216: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v217: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v218: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v219: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v220: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v221: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v222: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v223: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v224: OR2
        port map(Z0 => v119,
                 A0 => v117,
                 A1 => v120);
    
    v225: OR2
        port map(Z0 => v116,
                 A0 => v114,
                 A1 => v106);
    
    v226: OR2
        port map(Z0 => v113,
                 A0 => v110,
                 A1 => v111);
    
    v227: OR2
        port map(Z0 => v109,
                 A0 => v107,
                 A1 => v108);
    
    v228: AND3
        port map(Z0 => v105,
                 A0 => QI(0),
                 A1 => v121,
                 A2 => v122);
    
    v229: AND3
        port map(Z0 => v112,
                 A0 => QI(1),
                 A1 => v121,
                 A2 => v122);
    
    v230: AND3
        port map(Z0 => v115,
                 A0 => QI(2),
                 A1 => v121,
                 A2 => v122);
    
    v231: AND3
        port map(Z0 => v118,
                 A0 => QI(3),
                 A1 => v121,
                 A2 => v122);
    
    v232: FDC1
        port map(Q0 => QI(2),
                 D0 => v125,
                 CLK => CLK,
                 SD => SD);
    
    v233: FDC1
        port map(Q0 => QI(3),
                 D0 => v126,
                 CLK => CLK,
                 SD => SD);
    
    v234: AND3
        port map(Z0 => v107,
                 A0 => D0,
                 A1 => LD,
                 A2 => v122);
    
    v235: AND4
        port map(Z0 => v108,
                 A0 => v121,
                 A1 => CAI,
                 A2 => EN,
                 A3 => v122);
    
    v236: LXOR2
        port map(Z0 => v123,
                 A0 => v105,
                 A1 => v109);
    
    v237: LXOR2
        port map(Z0 => v124,
                 A0 => v112,
                 A1 => v113);
    
    v238: AND3
        port map(Z0 => v110,
                 A0 => D1,
                 A1 => LD,
                 A2 => v122);
    
    v239: INV
        port map(ZN0 => v121,
                 A0 => LD);
    
    v240: AND3
        port map(Z0 => v114,
                 A0 => D2,
                 A1 => LD,
                 A2 => v122);
    
    v241: LXOR2
        port map(Z0 => v125,
                 A0 => v115,
                 A1 => v116);
    
    v242: LXOR2
        port map(Z0 => v126,
                 A0 => v118,
                 A1 => v119);
    
    v243: AND3
        port map(Z0 => v117,
                 A0 => D3,
                 A1 => LD,
                 A2 => v122);
    
    v244: AND5
        port map(Z0 => v111,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v121,
                 A3 => EN,
                 A4 => v122);
    
    v245: AND8
        port map(Z0 => v132,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => v128,
                 A5 => CAI,
                 A6 => EN,
                 A7 => v141);
    
    v246: AND9
        port map(Z0 => v136,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => v128,
                 A6 => CAI,
                 A7 => EN,
                 A8 => v141);
    
    v247: AND10
        port map(Z0 => v137,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => v128,
                 A7 => CAI,
                 A8 => EN,
                 A9 => v141);
    
    v248: AND11
        port map(Z0 => v127,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => v128,
                 A8 => CAI,
                 A9 => EN,
                 A10 => v141);
    
    v249: INV
        port map(ZN0 => v141,
                 A0 => CS);
    
    v250: OR2
        port map(Z0 => v129,
                 A0 => v131,
                 A1 => v132);
    
    v251: OR2
        port map(Z0 => v133,
                 A0 => v135,
                 A1 => v136);
    
    v252: OR2
        port map(Z0 => v140,
                 A0 => v138,
                 A1 => v137);
    
    v253: OR2
        port map(Z0 => v142,
                 A0 => v144,
                 A1 => v127);
    
    v254: AND3
        port map(Z0 => v130,
                 A0 => QI(4),
                 A1 => v128,
                 A2 => v141);
    
    v255: AND3
        port map(Z0 => v134,
                 A0 => QI(5),
                 A1 => v128,
                 A2 => v141);
    
    v256: AND3
        port map(Z0 => v139,
                 A0 => QI(6),
                 A1 => v128,
                 A2 => v141);
    
    v257: AND3
        port map(Z0 => v143,
                 A0 => QI(7),
                 A1 => v128,
                 A2 => v141);
    
    v258: INV
        port map(ZN0 => v128,
                 A0 => LD);
    
    v259: LXOR2
        port map(Z0 => v145,
                 A0 => v130,
                 A1 => v129);
    
    v260: FDC1
        port map(Q0 => QI(4),
                 D0 => v145,
                 CLK => CLK,
                 SD => SD);
    
    v261: AND3
        port map(Z0 => v131,
                 A0 => D4,
                 A1 => LD,
                 A2 => v141);
    
    v262: LXOR2
        port map(Z0 => v146,
                 A0 => v134,
                 A1 => v133);
    
    v263: FDC1
        port map(Q0 => QI(5),
                 D0 => v146,
                 CLK => CLK,
                 SD => SD);
    
    v264: AND3
        port map(Z0 => v135,
                 A0 => D5,
                 A1 => LD,
                 A2 => v141);
    
    v265: AND3
        port map(Z0 => v138,
                 A0 => D6,
                 A1 => LD,
                 A2 => v141);
    
    v266: FDC1
        port map(Q0 => QI(6),
                 D0 => v147,
                 CLK => CLK,
                 SD => SD);
    
    v267: LXOR2
        port map(Z0 => v147,
                 A0 => v139,
                 A1 => v140);
    
    v268: LXOR2
        port map(Z0 => v148,
                 A0 => v143,
                 A1 => v142);
    
    v269: FDC1
        port map(Q0 => QI(7),
                 D0 => v148,
                 CLK => CLK,
                 SD => SD);
    
    v270: AND3
        port map(Z0 => v144,
                 A0 => D7,
                 A1 => LD,
                 A2 => v141);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUD4S is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         DNUP: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         CS: IN std_logic);
end CBUD4S;

architecture LATTICE_ARCH of CBUD4S is
    signal QI: std_logic_vector(0 to 3);
    signal v133: std_logic_vector(0 to 3);
    signal v111: std_logic;
    signal v106: std_logic;
    signal v124: std_logic;
    signal v104: std_logic;
    signal v120: std_logic;
    signal v105: std_logic;
    signal v119: std_logic;
    signal v121: std_logic;
    signal v114: std_logic;
    signal v107: std_logic;
    signal v128: std_logic;
    signal v113: std_logic;
    signal v108: std_logic;
    signal v123: std_logic;
    signal v112: std_logic;
    signal v110: std_logic;
    signal v125: std_logic;
    signal v122: std_logic;
    signal v118: std_logic;
    signal v109: std_logic;
    signal v127: std_logic;
    signal v116: std_logic;
    signal v126: std_logic;
    signal v117: std_logic;
    signal v100: std_logic;
    signal v102: std_logic;
    signal v103: std_logic;
    signal v101: std_logic;
    signal v115: std_logic;
    signal UP: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component OR3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : OR3 use entity LAT_VHD.OR3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
begin
    v177: FDE1
        port map(Q0 => QI(0),
                 D0 => v113,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v178: FDE1
        port map(Q0 => QI(1),
                 D0 => v114,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v179: OR2
        port map(Z0 => CAO,
                 A0 => v103,
                 A1 => v102);
    
    v180: INV
        port map(ZN0 => v101,
                 A0 => CS);
    
    v181: INV
        port map(ZN0 => UP,
                 A0 => DNUP);
    
    v182: AND7
        port map(Z0 => v102,
                 A0 => v133(0),
                 A1 => v133(1),
                 A2 => v133(2),
                 A3 => v133(3),
                 A4 => CAI,
                 A5 => EN,
                 A6 => DNUP);
    
    v183: AND7
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => CAI,
                 A5 => EN,
                 A6 => UP);
    
    v184: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v185: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v186: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v187: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v188: AND3
        port map(Z0 => v109,
                 A0 => QI(1),
                 A1 => v111,
                 A2 => v101);
    
    v189: AND3
        port map(Z0 => v100,
                 A0 => QI(0),
                 A1 => v111,
                 A2 => v101);
    
    v190: OR2
        port map(Z0 => v106,
                 A0 => v104,
                 A1 => v105);
    
    v191: OR3
        port map(Z0 => v110,
                 A0 => v107,
                 A1 => v108,
                 A2 => v112);
    
    v192: AND3
        port map(Z0 => v104,
                 A0 => D0,
                 A1 => LD,
                 A2 => v101);
    
    v193: AND4
        port map(Z0 => v105,
                 A0 => v111,
                 A1 => CAI,
                 A2 => EN,
                 A3 => v101);
    
    v194: LXOR2
        port map(Z0 => v113,
                 A0 => v100,
                 A1 => v106);
    
    v195: LXOR2
        port map(Z0 => v114,
                 A0 => v109,
                 A1 => v110);
    
    v196: AND3
        port map(Z0 => v107,
                 A0 => D1,
                 A1 => LD,
                 A2 => v101);
    
    v197: INV
        port map(ZN0 => v111,
                 A0 => LD);
    
    v198: AND6
        port map(Z0 => v108,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v111,
                 A3 => EN,
                 A4 => v101,
                 A5 => UP);
    
    v199: AND6
        port map(Z0 => v112,
                 A0 => v133(0),
                 A1 => CAI,
                 A2 => v111,
                 A3 => EN,
                 A4 => v101,
                 A5 => DNUP);
    
    v200: INV
        port map(ZN0 => v133(0),
                 A0 => QI(0));
    
    v201: INV
        port map(ZN0 => v133(1),
                 A0 => QI(1));
    
    v202: INV
        port map(ZN0 => v115,
                 A0 => CS);
    
    v203: AND3
        port map(Z0 => v117,
                 A0 => QI(2),
                 A1 => v124,
                 A2 => v115);
    
    v204: AND3
        port map(Z0 => v121,
                 A0 => QI(3),
                 A1 => v124,
                 A2 => v115);
    
    v205: OR3
        port map(Z0 => v118,
                 A0 => v116,
                 A1 => v119,
                 A2 => v125);
    
    v206: OR3
        port map(Z0 => v122,
                 A0 => v120,
                 A1 => v123,
                 A2 => v126);
    
    v207: FDE1
        port map(Q0 => QI(2),
                 D0 => v127,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v208: FDE1
        port map(Q0 => QI(3),
                 D0 => v128,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v209: INV
        port map(ZN0 => v124,
                 A0 => LD);
    
    v210: AND3
        port map(Z0 => v116,
                 A0 => D2,
                 A1 => LD,
                 A2 => v115);
    
    v211: LXOR2
        port map(Z0 => v127,
                 A0 => v117,
                 A1 => v118);
    
    v212: LXOR2
        port map(Z0 => v128,
                 A0 => v121,
                 A1 => v122);
    
    v213: AND3
        port map(Z0 => v120,
                 A0 => D3,
                 A1 => LD,
                 A2 => v115);
    
    v214: INV
        port map(ZN0 => v133(2),
                 A0 => QI(2));
    
    v215: INV
        port map(ZN0 => v133(3),
                 A0 => QI(3));
    
    v216: AND7
        port map(Z0 => v119,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => v124,
                 A3 => CAI,
                 A4 => EN,
                 A5 => v115,
                 A6 => UP);
    
    v217: AND7
        port map(Z0 => v125,
                 A0 => v133(0),
                 A1 => v133(1),
                 A2 => v124,
                 A3 => CAI,
                 A4 => EN,
                 A5 => v115,
                 A6 => DNUP);
    
    v218: AND8
        port map(Z0 => v123,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v124,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v115,
                 A7 => UP);
    
    v219: AND8
        port map(Z0 => v126,
                 A0 => v133(0),
                 A1 => v133(1),
                 A2 => v133(2),
                 A3 => v124,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v115,
                 A7 => DNUP);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CBUD8S is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         CAO: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         DNUP: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         CS: IN std_logic);
end CBUD8S;

architecture LATTICE_ARCH of CBUD8S is
    signal QI: std_logic_vector(0 to 7);
    signal v168: std_logic_vector(0 to 7);
    signal v114: std_logic;
    signal v109: std_logic;
    signal v127: std_logic;
    signal v133: std_logic;
    signal v107: std_logic;
    signal v146: std_logic;
    signal v123: std_logic;
    signal v108: std_logic;
    signal v137: std_logic;
    signal v122: std_logic;
    signal v124: std_logic;
    signal v117: std_logic;
    signal v110: std_logic;
    signal v131: std_logic;
    signal v116: std_logic;
    signal v111: std_logic;
    signal v151: std_logic;
    signal v134: std_logic;
    signal v126: std_logic;
    signal v115: std_logic;
    signal v113: std_logic;
    signal v158: std_logic;
    signal v152: std_logic;
    signal v147: std_logic;
    signal v138: std_logic;
    signal v128: std_logic;
    signal v125: std_logic;
    signal v121: std_logic;
    signal v112: std_logic;
    signal v139: std_logic;
    signal v130: std_logic;
    signal v144: std_logic;
    signal v143: std_logic;
    signal v140: std_logic;
    signal v135: std_logic;
    signal v119: std_logic;
    signal v150: std_logic;
    signal v136: std_logic;
    signal v159: std_logic;
    signal v155: std_logic;
    signal v142: std_logic;
    signal v129: std_logic;
    signal v156: std_logic;
    signal v120: std_logic;
    signal v153: std_logic;
    signal v148: std_logic;
    signal v145: std_logic;
    signal v154: std_logic;
    signal v149: std_logic;
    signal v141: std_logic;
    signal v157: std_logic;
    signal v103: std_logic;
    signal v105: std_logic;
    signal v132: std_logic;
    signal v106: std_logic;
    signal v104: std_logic;
    signal v118: std_logic;
    signal UP: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component AND11
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic);
    end component;
    for all : AND11 use entity LAT_VHD.AND11(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component OR3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : OR3 use entity LAT_VHD.OR3(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component LXOR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : LXOR2 use entity LAT_VHD.LXOR2(LATTICE_ARCH);
    
    component AND6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : AND6 use entity LAT_VHD.AND6(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component AND8
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic);
    end component;
    for all : AND8 use entity LAT_VHD.AND8(LATTICE_ARCH);
    
    component AND9
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic);
    end component;
    for all : AND9 use entity LAT_VHD.AND9(LATTICE_ARCH);
    
    component AND10
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic);
    end component;
    for all : AND10 use entity LAT_VHD.AND10(LATTICE_ARCH);
    
    component AND12
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic;
             A7: IN std_logic;
             A8: IN std_logic;
             A9: IN std_logic;
             A10: IN std_logic;
             A11: IN std_logic);
    end component;
    for all : AND12 use entity LAT_VHD.AND12(LATTICE_ARCH);
    
begin
    v252: FDE1
        port map(Q0 => QI(0),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v253: FDE1
        port map(Q0 => QI(1),
                 D0 => v117,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v254: OR2
        port map(Z0 => CAO,
                 A0 => v106,
                 A1 => v105);
    
    v255: AND11
        port map(Z0 => v106,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => QI(7),
                 A8 => CAI,
                 A9 => EN,
                 A10 => UP);
    
    v256: AND11
        port map(Z0 => v105,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v168(2),
                 A3 => v168(3),
                 A4 => v168(4),
                 A5 => v168(5),
                 A6 => v168(6),
                 A7 => v168(7),
                 A8 => CAI,
                 A9 => EN,
                 A10 => DNUP);
    
    v257: INV
        port map(ZN0 => v104,
                 A0 => CS);
    
    v258: INV
        port map(ZN0 => UP,
                 A0 => DNUP);
    
    v259: BUF
        port map(Z0 => Q7,
                 A0 => QI(7));
    
    v260: BUF
        port map(Z0 => Q6,
                 A0 => QI(6));
    
    v261: BUF
        port map(Z0 => Q5,
                 A0 => QI(5));
    
    v262: BUF
        port map(Z0 => Q4,
                 A0 => QI(4));
    
    v263: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v264: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v265: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v266: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v267: AND3
        port map(Z0 => v103,
                 A0 => QI(0),
                 A1 => v114,
                 A2 => v104);
    
    v268: AND3
        port map(Z0 => v112,
                 A0 => QI(1),
                 A1 => v114,
                 A2 => v104);
    
    v269: OR3
        port map(Z0 => v113,
                 A0 => v110,
                 A1 => v111,
                 A2 => v115);
    
    v270: OR2
        port map(Z0 => v109,
                 A0 => v107,
                 A1 => v108);
    
    v271: AND3
        port map(Z0 => v107,
                 A0 => D0,
                 A1 => LD,
                 A2 => v104);
    
    v272: AND4
        port map(Z0 => v108,
                 A0 => v114,
                 A1 => CAI,
                 A2 => EN,
                 A3 => v104);
    
    v273: LXOR2
        port map(Z0 => v116,
                 A0 => v103,
                 A1 => v109);
    
    v274: LXOR2
        port map(Z0 => v117,
                 A0 => v112,
                 A1 => v113);
    
    v275: AND3
        port map(Z0 => v110,
                 A0 => D1,
                 A1 => LD,
                 A2 => v104);
    
    v276: INV
        port map(ZN0 => v114,
                 A0 => LD);
    
    v277: AND6
        port map(Z0 => v111,
                 A0 => QI(0),
                 A1 => CAI,
                 A2 => v114,
                 A3 => EN,
                 A4 => v104,
                 A5 => UP);
    
    v278: AND6
        port map(Z0 => v115,
                 A0 => v168(0),
                 A1 => CAI,
                 A2 => v114,
                 A3 => EN,
                 A4 => v104,
                 A5 => DNUP);
    
    v279: INV
        port map(ZN0 => v168(0),
                 A0 => QI(0));
    
    v280: INV
        port map(ZN0 => v168(1),
                 A0 => QI(1));
    
    v281: INV
        port map(ZN0 => v118,
                 A0 => CS);
    
    v282: AND3
        port map(Z0 => v124,
                 A0 => QI(3),
                 A1 => v127,
                 A2 => v118);
    
    v283: AND3
        port map(Z0 => v120,
                 A0 => QI(2),
                 A1 => v127,
                 A2 => v118);
    
    v284: OR3
        port map(Z0 => v125,
                 A0 => v123,
                 A1 => v126,
                 A2 => v129);
    
    v285: OR3
        port map(Z0 => v121,
                 A0 => v119,
                 A1 => v122,
                 A2 => v128);
    
    v286: FDE1
        port map(Q0 => QI(2),
                 D0 => v130,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v287: FDE1
        port map(Q0 => QI(3),
                 D0 => v131,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v288: INV
        port map(ZN0 => v127,
                 A0 => LD);
    
    v289: AND3
        port map(Z0 => v119,
                 A0 => D2,
                 A1 => LD,
                 A2 => v118);
    
    v290: LXOR2
        port map(Z0 => v130,
                 A0 => v120,
                 A1 => v121);
    
    v291: LXOR2
        port map(Z0 => v131,
                 A0 => v124,
                 A1 => v125);
    
    v292: AND3
        port map(Z0 => v123,
                 A0 => D3,
                 A1 => LD,
                 A2 => v118);
    
    v293: INV
        port map(ZN0 => v168(2),
                 A0 => QI(2));
    
    v294: INV
        port map(ZN0 => v168(3),
                 A0 => QI(3));
    
    v295: AND7
        port map(Z0 => v122,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => v127,
                 A3 => CAI,
                 A4 => EN,
                 A5 => v118,
                 A6 => UP);
    
    v296: AND7
        port map(Z0 => v128,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v127,
                 A3 => CAI,
                 A4 => EN,
                 A5 => v118,
                 A6 => DNUP);
    
    v297: AND8
        port map(Z0 => v126,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => v127,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v118,
                 A7 => UP);
    
    v298: AND8
        port map(Z0 => v129,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v168(2),
                 A3 => v127,
                 A4 => CAI,
                 A5 => EN,
                 A6 => v118,
                 A7 => DNUP);
    
    v299: INV
        port map(ZN0 => v133,
                 A0 => LD);
    
    v300: INV
        port map(ZN0 => v134,
                 A0 => CS);
    
    v301: AND3
        port map(Z0 => v132,
                 A0 => QI(5),
                 A1 => v133,
                 A2 => v134);
    
    v302: AND3
        port map(Z0 => v137,
                 A0 => QI(4),
                 A1 => v133,
                 A2 => v134);
    
    v303: OR3
        port map(Z0 => v141,
                 A0 => v142,
                 A1 => v143,
                 A2 => v140);
    
    v304: OR3
        port map(Z0 => v136,
                 A0 => v138,
                 A1 => v139,
                 A2 => v135);
    
    v305: INV
        port map(ZN0 => v168(4),
                 A0 => QI(4));
    
    v306: LXOR2
        port map(Z0 => v144,
                 A0 => v137,
                 A1 => v136);
    
    v307: FDE1
        port map(Q0 => QI(4),
                 D0 => v144,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v308: AND3
        port map(Z0 => v138,
                 A0 => D4,
                 A1 => LD,
                 A2 => v134);
    
    v309: AND9
        port map(Z0 => v139,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => v133,
                 A5 => CAI,
                 A6 => EN,
                 A7 => v134,
                 A8 => UP);
    
    v310: AND9
        port map(Z0 => v135,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v168(2),
                 A3 => v168(3),
                 A4 => v133,
                 A5 => CAI,
                 A6 => EN,
                 A7 => v134,
                 A8 => DNUP);
    
    v311: INV
        port map(ZN0 => v168(5),
                 A0 => QI(5));
    
    v312: LXOR2
        port map(Z0 => v145,
                 A0 => v132,
                 A1 => v141);
    
    v313: FDE1
        port map(Q0 => QI(5),
                 D0 => v145,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v314: AND3
        port map(Z0 => v142,
                 A0 => D5,
                 A1 => LD,
                 A2 => v134);
    
    v315: AND10
        port map(Z0 => v143,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => v133,
                 A6 => CAI,
                 A7 => EN,
                 A8 => v134,
                 A9 => UP);
    
    v316: AND10
        port map(Z0 => v140,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v168(2),
                 A3 => v168(3),
                 A4 => v168(4),
                 A5 => v133,
                 A6 => CAI,
                 A7 => EN,
                 A8 => v134,
                 A9 => DNUP);
    
    v317: INV
        port map(ZN0 => v146,
                 A0 => LD);
    
    v318: INV
        port map(ZN0 => v147,
                 A0 => CS);
    
    v319: AND3
        port map(Z0 => v156,
                 A0 => QI(7),
                 A1 => v146,
                 A2 => v147);
    
    v320: AND3
        port map(Z0 => v151,
                 A0 => QI(6),
                 A1 => v146,
                 A2 => v147);
    
    v321: OR3
        port map(Z0 => v155,
                 A0 => v157,
                 A1 => v154,
                 A2 => v153);
    
    v322: OR3
        port map(Z0 => v152,
                 A0 => v150,
                 A1 => v149,
                 A2 => v148);
    
    v323: AND3
        port map(Z0 => v150,
                 A0 => D6,
                 A1 => LD,
                 A2 => v147);
    
    v324: FDE1
        port map(Q0 => QI(6),
                 D0 => v158,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v325: LXOR2
        port map(Z0 => v158,
                 A0 => v151,
                 A1 => v152);
    
    v326: INV
        port map(ZN0 => v168(6),
                 A0 => QI(6));
    
    v327: AND11
        port map(Z0 => v149,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => v146,
                 A7 => CAI,
                 A8 => EN,
                 A9 => v147,
                 A10 => UP);
    
    v328: AND11
        port map(Z0 => v148,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v168(2),
                 A3 => v168(3),
                 A4 => v168(4),
                 A5 => v168(5),
                 A6 => v146,
                 A7 => CAI,
                 A8 => EN,
                 A9 => v147,
                 A10 => DNUP);
    
    v329: INV
        port map(ZN0 => v168(7),
                 A0 => QI(7));
    
    v330: LXOR2
        port map(Z0 => v159,
                 A0 => v156,
                 A1 => v155);
    
    v331: FDE1
        port map(Q0 => QI(7),
                 D0 => v159,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v332: AND3
        port map(Z0 => v157,
                 A0 => D7,
                 A1 => LD,
                 A2 => v147);
    
    v333: AND12
        port map(Z0 => v154,
                 A0 => QI(0),
                 A1 => QI(1),
                 A2 => QI(2),
                 A3 => QI(3),
                 A4 => QI(4),
                 A5 => QI(5),
                 A6 => QI(6),
                 A7 => v146,
                 A8 => CAI,
                 A9 => EN,
                 A10 => v147,
                 A11 => UP);
    
    v334: AND12
        port map(Z0 => v153,
                 A0 => v168(0),
                 A1 => v168(1),
                 A2 => v168(2),
                 A3 => v168(3),
                 A4 => v168(4),
                 A5 => v168(5),
                 A6 => v168(6),
                 A7 => v146,
                 A8 => CAI,
                 A9 => EN,
                 A10 => v147,
                 A11 => DNUP);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CGD34 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic);
end CGD34;

architecture LATTICE_ARCH of CGD34 is
    signal v125: std_logic_vector(0 to 3);
    signal QI: std_logic_vector(0 to 3);
    signal v111: std_logic;
    signal v109: std_logic;
    signal v113: std_logic;
    signal v114: std_logic;
    signal v108: std_logic;
    signal v115: std_logic;
    signal v110: std_logic;
    signal LOAD0: std_logic;
    signal LOAD1: std_logic;
    signal LOAD2: std_logic;
    signal LOAD3: std_logic;
    signal HOLD0: std_logic;
    signal HOLD1: std_logic;
    signal HOLD2: std_logic;
    signal HOLD3: std_logic;
    signal v100: std_logic;
    signal v101: std_logic;
    signal v107: std_logic;
    signal v103: std_logic;
    signal v104: std_logic;
    signal v116: std_logic;
    signal v112: std_logic;
    signal v105: std_logic;
    signal v118: std_logic;
    signal v106: std_logic;
    signal v119: std_logic;
    signal v102: std_logic;
    signal v117: std_logic;
    signal v120: std_logic;
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : OR6 use entity LAT_VHD.OR6(LATTICE_ARCH);
    
    component OR5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : OR5 use entity LAT_VHD.OR5(LATTICE_ARCH);
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
begin
    v167: AND5
        port map(Z0 => v106,
                 A0 => QI(3),
                 A1 => v125(2),
                 A2 => QI(0),
                 A3 => v107,
                 A4 => EN);
    
    v168: AND3
        port map(Z0 => HOLD0,
                 A0 => QI(0),
                 A1 => v107,
                 A2 => v102);
    
    v169: AND2
        port map(Z0 => LOAD0,
                 A0 => D0,
                 A1 => LD);
    
    v170: AND5
        port map(Z0 => v100,
                 A0 => v125(3),
                 A1 => v125(2),
                 A2 => QI(1),
                 A3 => v107,
                 A4 => EN);
    
    v171: AND5
        port map(Z0 => v109,
                 A0 => v125(3),
                 A1 => QI(2),
                 A2 => v125(1),
                 A3 => v107,
                 A4 => EN);
    
    v172: AND5
        port map(Z0 => v101,
                 A0 => QI(3),
                 A1 => QI(2),
                 A2 => QI(1),
                 A3 => v107,
                 A4 => EN);
    
    v173: AND5
        port map(Z0 => v103,
                 A0 => QI(3),
                 A1 => v125(2),
                 A2 => v125(1),
                 A3 => v107,
                 A4 => EN);
    
    v174: AND3
        port map(Z0 => HOLD1,
                 A0 => QI(1),
                 A1 => v107,
                 A2 => v102);
    
    v175: AND2
        port map(Z0 => LOAD1,
                 A0 => D1,
                 A1 => LD);
    
    v176: AND5
        port map(Z0 => v104,
                 A0 => v125(3),
                 A1 => QI(2),
                 A2 => QI(0),
                 A3 => v107,
                 A4 => EN);
    
    v177: INV
        port map(ZN0 => v107,
                 A0 => LD);
    
    v178: INV
        port map(ZN0 => v102,
                 A0 => EN);
    
    v179: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v180: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v181: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v182: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v183: OR6
        port map(Z0 => v108,
                 A0 => HOLD0,
                 A1 => LOAD0,
                 A2 => v100,
                 A3 => v109,
                 A4 => v101,
                 A5 => v103);
    
    v184: OR5
        port map(Z0 => v110,
                 A0 => HOLD1,
                 A1 => LOAD1,
                 A2 => v105,
                 A3 => v104,
                 A4 => v106);
    
    v185: FDE1
        port map(Q0 => QI(0),
                 D0 => v108,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v186: FDE1
        port map(Q0 => QI(1),
                 D0 => v110,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v187: INV
        port map(ZN0 => v125(1),
                 A0 => QI(1));
    
    v188: INV
        port map(ZN0 => v125(0),
                 A0 => QI(0));
    
    v189: AND4
        port map(Z0 => v105,
                 A0 => QI(1),
                 A1 => v125(0),
                 A2 => v107,
                 A3 => EN);
    
    v190: INV
        port map(ZN0 => v118,
                 A0 => LD);
    
    v191: INV
        port map(ZN0 => v117,
                 A0 => EN);
    
    v192: OR5
        port map(Z0 => v116,
                 A0 => HOLD2,
                 A1 => LOAD2,
                 A2 => v115,
                 A3 => v114,
                 A4 => v113);
    
    v193: OR5
        port map(Z0 => v112,
                 A0 => HOLD3,
                 A1 => LOAD3,
                 A2 => v111,
                 A3 => v119,
                 A4 => v120);
    
    v194: INV
        port map(ZN0 => v125(3),
                 A0 => QI(3));
    
    v195: AND5
        port map(Z0 => v115,
                 A0 => QI(3),
                 A1 => QI(1),
                 A2 => v125(0),
                 A3 => v118,
                 A4 => EN);
    
    v196: AND2
        port map(Z0 => LOAD2,
                 A0 => D2,
                 A1 => LD);
    
    v197: INV
        port map(ZN0 => v125(2),
                 A0 => QI(2));
    
    v198: AND4
        port map(Z0 => v114,
                 A0 => QI(2),
                 A1 => v125(1),
                 A2 => v118,
                 A3 => EN);
    
    v199: AND3
        port map(Z0 => HOLD3,
                 A0 => QI(3),
                 A1 => v118,
                 A2 => v117);
    
    v200: AND2
        port map(Z0 => LOAD3,
                 A0 => D3,
                 A1 => LD);
    
    v201: AND5
        port map(Z0 => v111,
                 A0 => v125(2),
                 A1 => v125(1),
                 A2 => v125(0),
                 A3 => v118,
                 A4 => EN);
    
    v202: AND4
        port map(Z0 => v119,
                 A0 => QI(3),
                 A1 => QI(0),
                 A2 => v118,
                 A3 => EN);
    
    v203: AND4
        port map(Z0 => v120,
                 A0 => QI(3),
                 A1 => QI(1),
                 A2 => v118,
                 A3 => EN);
    
    v204: AND4
        port map(Z0 => v113,
                 A0 => QI(2),
                 A1 => QI(0),
                 A2 => v118,
                 A3 => EN);
    
    v205: AND3
        port map(Z0 => HOLD2,
                 A0 => QI(2),
                 A1 => v118,
                 A2 => v117);
    
    v206: FDE1
        port map(Q0 => QI(2),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v207: FDE1
        port map(Q0 => QI(3),
                 D0 => v112,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CGU34 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic);
end CGU34;

architecture LATTICE_ARCH of CGU34 is
    signal QI: std_logic_vector(0 to 3);
    signal v125: std_logic_vector(0 to 3);
    signal v111: std_logic;
    signal v109: std_logic;
    signal v113: std_logic;
    signal v114: std_logic;
    signal v108: std_logic;
    signal v115: std_logic;
    signal v110: std_logic;
    signal LOAD0: std_logic;
    signal LOAD1: std_logic;
    signal LOAD2: std_logic;
    signal LOAD3: std_logic;
    signal HOLD0: std_logic;
    signal HOLD1: std_logic;
    signal HOLD2: std_logic;
    signal HOLD3: std_logic;
    signal v100: std_logic;
    signal v101: std_logic;
    signal v107: std_logic;
    signal v103: std_logic;
    signal v104: std_logic;
    signal v116: std_logic;
    signal v112: std_logic;
    signal v105: std_logic;
    signal v118: std_logic;
    signal v106: std_logic;
    signal v119: std_logic;
    signal v102: std_logic;
    signal v117: std_logic;
    signal v120: std_logic;
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : OR6 use entity LAT_VHD.OR6(LATTICE_ARCH);
    
    component OR5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : OR5 use entity LAT_VHD.OR5(LATTICE_ARCH);
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
begin
    v167: AND5
        port map(Z0 => v106,
                 A0 => QI(3),
                 A1 => QI(2),
                 A2 => QI(0),
                 A3 => v107,
                 A4 => EN);
    
    v168: AND3
        port map(Z0 => HOLD0,
                 A0 => QI(0),
                 A1 => v107,
                 A2 => v102);
    
    v169: AND2
        port map(Z0 => LOAD0,
                 A0 => D0,
                 A1 => LD);
    
    v170: AND5
        port map(Z0 => v100,
                 A0 => v125(3),
                 A1 => v125(2),
                 A2 => v125(1),
                 A3 => v107,
                 A4 => EN);
    
    v171: AND5
        port map(Z0 => v109,
                 A0 => v125(3),
                 A1 => QI(2),
                 A2 => QI(1),
                 A3 => v107,
                 A4 => EN);
    
    v172: AND5
        port map(Z0 => v101,
                 A0 => QI(3),
                 A1 => QI(2),
                 A2 => v125(1),
                 A3 => v107,
                 A4 => EN);
    
    v173: AND5
        port map(Z0 => v103,
                 A0 => QI(3),
                 A1 => v125(2),
                 A2 => QI(1),
                 A3 => v107,
                 A4 => EN);
    
    v174: AND3
        port map(Z0 => HOLD1,
                 A0 => QI(1),
                 A1 => v107,
                 A2 => v102);
    
    v175: AND2
        port map(Z0 => LOAD1,
                 A0 => D1,
                 A1 => LD);
    
    v176: AND5
        port map(Z0 => v104,
                 A0 => v125(3),
                 A1 => v125(2),
                 A2 => QI(0),
                 A3 => v107,
                 A4 => EN);
    
    v177: INV
        port map(ZN0 => v107,
                 A0 => LD);
    
    v178: INV
        port map(ZN0 => v102,
                 A0 => EN);
    
    v179: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v180: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v181: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v182: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v183: OR6
        port map(Z0 => v108,
                 A0 => HOLD0,
                 A1 => LOAD0,
                 A2 => v100,
                 A3 => v109,
                 A4 => v101,
                 A5 => v103);
    
    v184: OR5
        port map(Z0 => v110,
                 A0 => HOLD1,
                 A1 => LOAD1,
                 A2 => v105,
                 A3 => v104,
                 A4 => v106);
    
    v185: FDE1
        port map(Q0 => QI(0),
                 D0 => v108,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v186: FDE1
        port map(Q0 => QI(1),
                 D0 => v110,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v187: INV
        port map(ZN0 => v125(1),
                 A0 => QI(1));
    
    v188: INV
        port map(ZN0 => v125(0),
                 A0 => QI(0));
    
    v189: AND4
        port map(Z0 => v105,
                 A0 => QI(1),
                 A1 => v125(0),
                 A2 => v107,
                 A3 => EN);
    
    v190: INV
        port map(ZN0 => v118,
                 A0 => LD);
    
    v191: INV
        port map(ZN0 => v117,
                 A0 => EN);
    
    v192: OR5
        port map(Z0 => v112,
                 A0 => HOLD3,
                 A1 => LOAD3,
                 A2 => v111,
                 A3 => v119,
                 A4 => v120);
    
    v193: OR5
        port map(Z0 => v116,
                 A0 => HOLD2,
                 A1 => LOAD2,
                 A2 => v115,
                 A3 => v114,
                 A4 => v113);
    
    v194: INV
        port map(ZN0 => v125(3),
                 A0 => QI(3));
    
    v195: AND5
        port map(Z0 => v115,
                 A0 => v125(3),
                 A1 => QI(1),
                 A2 => v125(0),
                 A3 => v118,
                 A4 => EN);
    
    v196: AND2
        port map(Z0 => LOAD2,
                 A0 => D2,
                 A1 => LD);
    
    v197: INV
        port map(ZN0 => v125(2),
                 A0 => QI(2));
    
    v198: AND4
        port map(Z0 => v114,
                 A0 => QI(2),
                 A1 => v125(1),
                 A2 => v118,
                 A3 => EN);
    
    v199: AND3
        port map(Z0 => HOLD3,
                 A0 => QI(3),
                 A1 => v118,
                 A2 => v117);
    
    v200: AND2
        port map(Z0 => LOAD3,
                 A0 => D3,
                 A1 => LD);
    
    v201: AND5
        port map(Z0 => v111,
                 A0 => QI(2),
                 A1 => v125(1),
                 A2 => v125(0),
                 A3 => v118,
                 A4 => EN);
    
    v202: AND4
        port map(Z0 => v119,
                 A0 => QI(3),
                 A1 => QI(0),
                 A2 => v118,
                 A3 => EN);
    
    v203: AND4
        port map(Z0 => v120,
                 A0 => QI(3),
                 A1 => QI(1),
                 A2 => v118,
                 A3 => EN);
    
    v204: AND4
        port map(Z0 => v113,
                 A0 => QI(2),
                 A1 => QI(0),
                 A2 => v118,
                 A3 => EN);
    
    v205: AND3
        port map(Z0 => HOLD2,
                 A0 => QI(2),
                 A1 => v118,
                 A2 => v117);
    
    v206: FDE1
        port map(Q0 => QI(2),
                 D0 => v116,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v207: FDE1
        port map(Q0 => QI(3),
                 D0 => v112,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity CGUD4S is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         DNUP: IN std_logic;
         CD: IN std_logic;
         CS: IN std_logic);
end CGUD4S;

architecture LATTICE_ARCH of CGUD4S is
    signal v145: std_logic_vector(0 to 3);
    signal QI: std_logic_vector(0 to 3);
    signal v129: std_logic;
    signal v114: std_logic;
    signal v127: std_logic;
    signal v135: std_logic;
    signal v130: std_logic;
    signal v136: std_logic;
    signal v134: std_logic;
    signal v131: std_logic;
    signal v137: std_logic;
    signal v133: std_logic;
    signal v128: std_logic;
    signal v118: std_logic;
    signal v132: std_logic;
    signal v122: std_logic;
    signal LOAD0: std_logic;
    signal LOAD1: std_logic;
    signal LOAD2: std_logic;
    signal LOAD3: std_logic;
    signal HOLD0: std_logic;
    signal HOLD1: std_logic;
    signal HOLD2: std_logic;
    signal HOLD3: std_logic;
    signal v100: std_logic;
    signal v102: std_logic;
    signal v116: std_logic;
    signal v107: std_logic;
    signal v117: std_logic;
    signal v108: std_logic;
    signal v112: std_logic;
    signal v103: std_logic;
    signal v109: std_logic;
    signal v138: std_logic;
    signal v113: std_logic;
    signal v104: std_logic;
    signal v115: std_logic;
    signal v105: std_logic;
    signal v140: std_logic;
    signal v110: std_logic;
    signal v106: std_logic;
    signal v111: std_logic;
    signal v101: std_logic;
    signal v123: std_logic;
    signal v139: std_logic;
    signal v124: std_logic;
    signal v119: std_logic;
    signal v120: std_logic;
    signal v125: std_logic;
    signal v121: std_logic;
    signal v126: std_logic;
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component AND7
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic;
             A6: IN std_logic);
    end component;
    for all : AND7 use entity LAT_VHD.AND7(LATTICE_ARCH);
    
    component OR4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all : OR4 use entity LAT_VHD.OR4(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component OR6
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic;
             A5: IN std_logic);
    end component;
    for all : OR6 use entity LAT_VHD.OR6(LATTICE_ARCH);
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component OR3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all : OR3 use entity LAT_VHD.OR3(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all : AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
begin
    v207: INV
        port map(ZN0 => v101,
                 A0 => EN);
    
    v208: AND4
        port map(Z0 => HOLD0,
                 A0 => QI(0),
                 A1 => v102,
                 A2 => v101,
                 A3 => v105);
    
    v209: AND3
        port map(Z0 => LOAD0,
                 A0 => D0,
                 A1 => LD,
                 A2 => v105);
    
    v210: AND7
        port map(Z0 => v100,
                 A0 => v145(3),
                 A1 => v145(2),
                 A2 => v145(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => v113);
    
    v211: AND7
        port map(Z0 => v114,
                 A0 => v145(3),
                 A1 => QI(2),
                 A2 => QI(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => v113);
    
    v212: AND7
        port map(Z0 => v103,
                 A0 => QI(3),
                 A1 => QI(2),
                 A2 => v145(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => v113);
    
    v213: AND7
        port map(Z0 => v104,
                 A0 => QI(3),
                 A1 => v145(2),
                 A2 => QI(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => v113);
    
    v214: INV
        port map(ZN0 => v102,
                 A0 => LD);
    
    v215: INV
        port map(ZN0 => v105,
                 A0 => CS);
    
    v216: AND7
        port map(Z0 => v109,
                 A0 => v145(3),
                 A1 => v145(2),
                 A2 => QI(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => DNUP);
    
    v217: AND7
        port map(Z0 => v107,
                 A0 => v145(3),
                 A1 => QI(2),
                 A2 => v145(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => DNUP);
    
    v218: AND7
        port map(Z0 => v106,
                 A0 => QI(3),
                 A1 => QI(2),
                 A2 => QI(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => DNUP);
    
    v219: AND7
        port map(Z0 => v108,
                 A0 => QI(3),
                 A1 => v145(2),
                 A2 => v145(1),
                 A3 => v102,
                 A4 => EN,
                 A5 => v105,
                 A6 => DNUP);
    
    v220: OR4
        port map(Z0 => v111,
                 A0 => v109,
                 A1 => v107,
                 A2 => v106,
                 A3 => v108);
    
    v221: OR2
        port map(Z0 => v112,
                 A0 => v110,
                 A1 => v111);
    
    v222: INV
        port map(ZN0 => v113,
                 A0 => DNUP);
    
    v223: BUF
        port map(Z0 => Q3,
                 A0 => QI(3));
    
    v224: BUF
        port map(Z0 => Q2,
                 A0 => QI(2));
    
    v225: BUF
        port map(Z0 => Q1,
                 A0 => QI(1));
    
    v226: BUF
        port map(Z0 => Q0,
                 A0 => QI(0));
    
    v227: OR6
        port map(Z0 => v110,
                 A0 => HOLD0,
                 A1 => LOAD0,
                 A2 => v100,
                 A3 => v114,
                 A4 => v103,
                 A5 => v104);
    
    v228: FDE1
        port map(Q0 => QI(0),
                 D0 => v112,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v229: INV
        port map(ZN0 => v145(0),
                 A0 => QI(0));
    
    v230: INV
        port map(ZN0 => v126,
                 A0 => DNUP);
    
    v231: FDE1
        port map(Q0 => QI(1),
                 D0 => v125,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v232: OR3
        port map(Z0 => v123,
                 A0 => HOLD1,
                 A1 => LOAD1,
                 A2 => v117);
    
    v233: INV
        port map(ZN0 => v145(1),
                 A0 => QI(1));
    
    v234: AND5
        port map(Z0 => v117,
                 A0 => QI(1),
                 A1 => v145(0),
                 A2 => v115,
                 A3 => EN,
                 A4 => v118);
    
    v235: AND4
        port map(Z0 => HOLD1,
                 A0 => QI(1),
                 A1 => v115,
                 A2 => v122,
                 A3 => v118);
    
    v236: INV
        port map(ZN0 => v122,
                 A0 => EN);
    
    v237: AND3
        port map(Z0 => LOAD1,
                 A0 => D1,
                 A1 => LD,
                 A2 => v118);
    
    v238: INV
        port map(ZN0 => v118,
                 A0 => CS);
    
    v239: INV
        port map(ZN0 => v115,
                 A0 => LD);
    
    v240: AND7
        port map(Z0 => v116,
                 A0 => v145(3),
                 A1 => v145(2),
                 A2 => QI(0),
                 A3 => v115,
                 A4 => EN,
                 A5 => v118,
                 A6 => v126);
    
    v241: AND7
        port map(Z0 => v119,
                 A0 => QI(3),
                 A1 => QI(2),
                 A2 => QI(0),
                 A3 => v115,
                 A4 => EN,
                 A5 => v118,
                 A6 => v126);
    
    v242: AND7
        port map(Z0 => v120,
                 A0 => v145(3),
                 A1 => QI(2),
                 A2 => QI(0),
                 A3 => v115,
                 A4 => EN,
                 A5 => v118,
                 A6 => DNUP);
    
    v243: AND7
        port map(Z0 => v121,
                 A0 => QI(3),
                 A1 => v145(2),
                 A2 => QI(0),
                 A3 => v115,
                 A4 => EN,
                 A5 => v118,
                 A6 => DNUP);
    
    v244: OR4
        port map(Z0 => v124,
                 A0 => v116,
                 A1 => v119,
                 A2 => v120,
                 A3 => v121);
    
    v245: OR2
        port map(Z0 => v125,
                 A0 => v123,
                 A1 => v124);
    
    v246: INV
        port map(ZN0 => v139,
                 A0 => EN);
    
    v247: AND4
        port map(Z0 => HOLD2,
                 A0 => QI(2),
                 A1 => v140,
                 A2 => v139,
                 A3 => v127);
    
    v248: AND3
        port map(Z0 => LOAD2,
                 A0 => D2,
                 A1 => LD,
                 A2 => v127);
    
    v249: AND5
        port map(Z0 => v136,
                 A0 => QI(2),
                 A1 => v145(1),
                 A2 => v140,
                 A3 => EN,
                 A4 => v127);
    
    v250: AND5
        port map(Z0 => v135,
                 A0 => QI(2),
                 A1 => QI(0),
                 A2 => v140,
                 A3 => EN,
                 A4 => v127);
    
    v251: AND7
        port map(Z0 => v137,
                 A0 => v145(3),
                 A1 => QI(1),
                 A2 => v145(0),
                 A3 => v140,
                 A4 => EN,
                 A5 => v127,
                 A6 => v129);
    
    v252: AND7
        port map(Z0 => v128,
                 A0 => QI(3),
                 A1 => QI(1),
                 A2 => v145(0),
                 A3 => v140,
                 A4 => EN,
                 A5 => v127,
                 A6 => DNUP);
    
    v253: AND4
        port map(Z0 => HOLD3,
                 A0 => QI(3),
                 A1 => v140,
                 A2 => v139,
                 A3 => v127);
    
    v254: AND7
        port map(Z0 => v134,
                 A0 => v145(2),
                 A1 => v145(1),
                 A2 => v145(0),
                 A3 => v140,
                 A4 => EN,
                 A5 => v127,
                 A6 => DNUP);
    
    v255: INV
        port map(ZN0 => v127,
                 A0 => CS);
    
    v256: AND7
        port map(Z0 => v132,
                 A0 => QI(2),
                 A1 => v145(1),
                 A2 => v145(0),
                 A3 => v140,
                 A4 => EN,
                 A5 => v127,
                 A6 => v129);
    
    v257: AND5
        port map(Z0 => v131,
                 A0 => QI(3),
                 A1 => QI(0),
                 A2 => v140,
                 A3 => EN,
                 A4 => v127);
    
    v258: INV
        port map(ZN0 => v140,
                 A0 => LD);
    
    v259: AND5
        port map(Z0 => v130,
                 A0 => QI(3),
                 A1 => QI(1),
                 A2 => v140,
                 A3 => EN,
                 A4 => v127);
    
    v260: AND3
        port map(Z0 => LOAD3,
                 A0 => D3,
                 A1 => LD,
                 A2 => v127);
    
    v261: INV
        port map(ZN0 => v145(3),
                 A0 => QI(3));
    
    v262: FDE1
        port map(Q0 => QI(3),
                 D0 => v133,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v263: INV
        port map(ZN0 => v129,
                 A0 => DNUP);
    
    v264: OR6
        port map(Z0 => v133,
                 A0 => HOLD3,
                 A1 => LOAD3,
                 A2 => v132,
                 A3 => v134,
                 A4 => v131,
                 A5 => v130);
    
    v265: OR6
        port map(Z0 => v138,
                 A0 => HOLD2,
                 A1 => LOAD2,
                 A2 => v137,
                 A3 => v128,
                 A4 => v136,
                 A5 => v135);
    
    v266: INV
        port map(ZN0 => v145(2),
                 A0 => QI(2));
    
    v267: FDE1
        port map(Q0 => QI(2),
                 D0 => v138,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FD14E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FD14E;

architecture LATTICE_ARCH of FD14E is
    
    component FD11E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: FD11E use entity LAT_VHD.FD11E(LATTICE_ARCH);
    
begin
    v110: FD11E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN);
    
    v111: FD11E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 EN => EN);
    
    v112: FD11E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 EN => EN);
    
    v113: FD11E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FD18E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FD18E;

architecture LATTICE_ARCH of FD18E is
    
    component FD11E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: FD11E use entity LAT_VHD.FD11E(LATTICE_ARCH);
    
begin
    v114: FD11E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN);
    
    v115: FD11E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 EN => EN);
    
    v116: FD11E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 EN => EN);
    
    v117: FD11E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 EN => EN);
    
    v118: FD11E
        port map(Q0 => Q7,
                 D0 => D7,
                 CLK => CLK,
                 EN => EN);
    
    v119: FD11E
        port map(Q0 => Q6,
                 D0 => D6,
                 CLK => CLK,
                 EN => EN);
    
    v120: FD11E
        port map(Q0 => Q5,
                 D0 => D5,
                 CLK => CLK,
                 EN => EN);
    
    v121: FD11E
        port map(Q0 => Q4,
                 D0 => D4,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FD24E is
    port(CD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FD24E;

architecture LATTICE_ARCH of FD24E is
    
    component FD21E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FD21E use entity LAT_VHD.FD21E(LATTICE_ARCH);
    
begin
    v111: FD21E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v112: FD21E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v113: FD21E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v114: FD21E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FD28E is
    port(CD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FD28E;

architecture LATTICE_ARCH of FD28E is
    
    component FD21E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FD21E use entity LAT_VHD.FD21E(LATTICE_ARCH);
    
begin
    v115: FD21E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v116: FD21E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v117: FD21E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v118: FD21E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v119: FD21E
        port map(Q0 => Q4,
                 D0 => D4,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v120: FD21E
        port map(Q0 => Q5,
                 D0 => D5,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v121: FD21E
        port map(Q0 => Q6,
                 D0 => D6,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    v122: FD21E
        port map(Q0 => Q7,
                 D0 => D7,
                 CLK => CLK,
                 EN => EN,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDC4 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic);
end FDC4;

architecture LATTICE_ARCH of FDC4 is
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
begin
    v107: FDC1
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD);
    
    v108: FDC1
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD);
    
    v109: FDC1
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD);
    
    v110: FDC1
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDC4E is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FDC4E;

architecture LATTICE_ARCH of FDC4E is
    
    component FDC1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : FDC1E use entity LAT_VHD.FDC1E(LATTICE_ARCH);
    
begin
    v111: FDC1E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v112: FDC1E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v113: FDC1E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v114: FDC1E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDC8 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CLK: IN std_logic);
end FDC8;

architecture LATTICE_ARCH of FDC8 is
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
begin
    v111: FDC1
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD);
    
    v112: FDC1
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD);
    
    v113: FDC1
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD);
    
    v114: FDC1
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD);
    
    v115: FDC1
        port map(Q0 => Q4,
                 D0 => D4,
                 CLK => CLK,
                 SD => SD);
    
    v116: FDC1
        port map(Q0 => Q5,
                 D0 => D5,
                 CLK => CLK,
                 SD => SD);
    
    v117: FDC1
        port map(Q0 => Q6,
                 D0 => D6,
                 CLK => CLK,
                 SD => SD);
    
    v118: FDC1
        port map(Q0 => Q7,
                 D0 => D7,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDC8E is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FDC8E;

architecture LATTICE_ARCH of FDC8E is
    
    component FDC1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : FDC1E use entity LAT_VHD.FDC1E(LATTICE_ARCH);
    
begin
    v115: FDC1E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v116: FDC1E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v117: FDC1E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v118: FDC1E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v119: FDC1E
        port map(Q0 => Q7,
                 D0 => D7,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v120: FDC1E
        port map(Q0 => Q6,
                 D0 => D6,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v121: FDC1E
        port map(Q0 => Q5,
                 D0 => D5,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    v122: FDC1E
        port map(Q0 => Q4,
                 D0 => D4,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDE4 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic);
end FDE4;

architecture LATTICE_ARCH of FDE4 is
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
begin
    v104: FDE1
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v105: FDE1
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v106: FDE1
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v107: FDE1
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDE4E is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FDE4E;

architecture LATTICE_ARCH of FDE4E is
    
    component FDE1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : FDE1E use entity LAT_VHD.FDE1E(LATTICE_ARCH);
    
begin
    v108: FDE1E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v109: FDE1E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v110: FDE1E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v111: FDE1E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDE8 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CLK: IN std_logic);
end FDE8;

architecture LATTICE_ARCH of FDE8 is
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
begin
    v108: FDE1
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v109: FDE1
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v110: FDE1
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v111: FDE1
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v112: FDE1
        port map(Q0 => Q4,
                 D0 => D4,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v113: FDE1
        port map(Q0 => Q5,
                 D0 => D5,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v114: FDE1
        port map(Q0 => Q6,
                 D0 => D6,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v115: FDE1
        port map(Q0 => Q7,
                 D0 => D7,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FDE8E is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         EN: IN std_logic;
         CLK: IN std_logic);
end FDE8E;

architecture LATTICE_ARCH of FDE8E is
    
    component FDE1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : FDE1E use entity LAT_VHD.FDE1E(LATTICE_ARCH);
    
begin
    v112: FDE1E
        port map(Q0 => Q3,
                 D0 => D3,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v113: FDE1E
        port map(Q0 => Q0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v114: FDE1E
        port map(Q0 => Q1,
                 D0 => D1,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v115: FDE1E
        port map(Q0 => Q2,
                 D0 => D2,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v116: FDE1E
        port map(Q0 => Q7,
                 D0 => D7,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v117: FDE1E
        port map(Q0 => Q6,
                 D0 => D6,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v118: FDE1E
        port map(Q0 => Q5,
                 D0 => D5,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v119: FDE1E
        port map(Q0 => Q4,
                 D0 => D4,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK61 is
    port(Q0: OUT std_logic;
         J0: IN std_logic;
         K0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic);
end FJK61;

architecture LATTICE_ARCH of FJK61 is
    signal v107: std_logic;
    signal v105: std_logic;
    signal v103: std_logic;
    signal v106: std_logic;
    signal v104: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);
    
    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
begin
    v114: FDC1
        port map(Q0 => v106,
                 D0 => v107,
                 CLK => CLK,
                 SD => SD);
    
    v115: NAND2
        port map(ZN0 => v103,
                 A0 => v105,
                 A1 => J0);
    
    v116: OR2
        port map(Z0 => v104,
                 A0 => v105,
                 A1 => K0);
    
    v117: NAND2
        port map(ZN0 => v107,
                 A0 => v103,
                 A1 => v104);
    
    v118: INV
        port map(ZN0 => v105,
                 A0 => v106);
    
    v119: BUF
        port map(Z0 => Q0,
                 A0 => v106);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK64 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         J0: IN std_logic;
         J1: IN std_logic;
         J2: IN std_logic;
         J3: IN std_logic;
         K0: IN std_logic;
         K1: IN std_logic;
         K2: IN std_logic;
         K3: IN std_logic;
         CLK: IN std_logic);
end FJK64;

architecture LATTICE_ARCH of FJK64 is
    signal v103,v104,v105,v106,v107: std_logic;
    signal v113,v114,v115,v116,v117: std_logic;
    signal v123,v124,v125,v126,v127: std_logic;
    signal v133,v134,v135,v136,v137: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);

    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);
 
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);

    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

begin
    vv101: FDC1 port map(Q0 => v106, D0 => v107, CLK => CLK, SD => SD);
    vv102: FDC1 port map(Q0 => v116, D0 => v117, CLK => CLK, SD => SD);
    vv103: FDC1 port map(Q0 => v126, D0 => v127, CLK => CLK, SD => SD);
    vv104: FDC1 port map(Q0 => v136, D0 => v137, CLK => CLK, SD => SD);

    vv105: NAND2 port map(ZN0 => v103, A0 => v105, A1 => J0);
    vv106: NAND2 port map(ZN0 => v113, A0 => v115, A1 => J1);
    vv107: NAND2 port map(ZN0 => v123, A0 => v125, A1 => J2);
    vv108: NAND2 port map(ZN0 => v133, A0 => v135, A1 => J3);
    
    vv109: OR2 port map(Z0 => v104, A0 => v105, A1 => K0);
    vv110: OR2 port map(Z0 => v114, A0 => v115, A1 => K1);
    vv111: OR2 port map(Z0 => v124, A0 => v125, A1 => K2);
    vv112: OR2 port map(Z0 => v134, A0 => v135, A1 => K3);

    vv113: NAND2 port map(ZN0 => v107, A0 => v103, A1 => v104);
    vv114: NAND2 port map(ZN0 => v117, A0 => v113, A1 => v114);
    vv115: NAND2 port map(ZN0 => v127, A0 => v123, A1 => v124);
    vv116: NAND2 port map(ZN0 => v137, A0 => v133, A1 => v134);

    vv117: INV port map(ZN0 => v105, A0 => v106);
    vv118: INV port map(ZN0 => v115, A0 => v116);
    vv119: INV port map(ZN0 => v125, A0 => v126);
    vv120: INV port map(ZN0 => v135, A0 => v136);

    vv121: BUF port map(Z0 => Q0, A0 => v106);
    vv122: BUF port map(Z0 => Q1, A0 => v116);
    vv123: BUF port map(Z0 => Q2, A0 => v126);
    vv124: BUF port map(Z0 => Q3, A0 => v136);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK68 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         J0: IN std_logic;
         J1: IN std_logic;
         J2: IN std_logic;
         J3: IN std_logic;
         J4: IN std_logic;
         J5: IN std_logic;
         J6: IN std_logic;
         J7: IN std_logic;
         K0: IN std_logic;
         K1: IN std_logic;
         K2: IN std_logic;
         K3: IN std_logic;
         K4: IN std_logic;
         K5: IN std_logic;
         K6: IN std_logic;
         K7: IN std_logic;
         CLK: IN std_logic);
end FJK68;

architecture LATTICE_ARCH of FJK68 is
    signal v103,v104,v105,v106,v107: std_logic;
    signal v113,v114,v115,v116,v117: std_logic;
    signal v123,v124,v125,v126,v127: std_logic;
    signal v133,v134,v135,v136,v137: std_logic;
    signal v143,v144,v145,v146,v147: std_logic;
    signal v153,v154,v155,v156,v157: std_logic;
    signal v163,v164,v165,v166,v167: std_logic;
    signal v173,v174,v175,v176,v177: std_logic;
    
    component FDC1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : FDC1 use entity LAT_VHD.FDC1(LATTICE_ARCH);

    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);
 
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);

    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

begin
    vv101: FDC1 port map(Q0 => v106, D0 => v107, CLK => CLK, SD => SD);
    vv102: FDC1 port map(Q0 => v116, D0 => v117, CLK => CLK, SD => SD);
    vv103: FDC1 port map(Q0 => v126, D0 => v127, CLK => CLK, SD => SD);
    vv104: FDC1 port map(Q0 => v136, D0 => v137, CLK => CLK, SD => SD);
    vv105: FDC1 port map(Q0 => v146, D0 => v147, CLK => CLK, SD => SD);
    vv106: FDC1 port map(Q0 => v156, D0 => v157, CLK => CLK, SD => SD);
    vv107: FDC1 port map(Q0 => v166, D0 => v167, CLK => CLK, SD => SD);
    vv108: FDC1 port map(Q0 => v176, D0 => v177, CLK => CLK, SD => SD);

    vv109: NAND2 port map(ZN0 => v103, A0 => v105, A1 => J0);
    vv110: NAND2 port map(ZN0 => v113, A0 => v115, A1 => J1);
    vv111: NAND2 port map(ZN0 => v123, A0 => v125, A1 => J2);
    vv112: NAND2 port map(ZN0 => v133, A0 => v135, A1 => J3);
    vv113: NAND2 port map(ZN0 => v143, A0 => v145, A1 => J4);
    vv114: NAND2 port map(ZN0 => v153, A0 => v155, A1 => J5);
    vv115: NAND2 port map(ZN0 => v163, A0 => v165, A1 => J6);
    vv116: NAND2 port map(ZN0 => v173, A0 => v175, A1 => J7);
    
    vv117: OR2 port map(Z0 => v104, A0 => v105, A1 => K0);
    vv118: OR2 port map(Z0 => v114, A0 => v115, A1 => K1);
    vv119: OR2 port map(Z0 => v124, A0 => v125, A1 => K2);
    vv120: OR2 port map(Z0 => v134, A0 => v135, A1 => K3);
    vv121: OR2 port map(Z0 => v144, A0 => v145, A1 => K4);
    vv122: OR2 port map(Z0 => v154, A0 => v155, A1 => K5);
    vv123: OR2 port map(Z0 => v164, A0 => v165, A1 => K6);
    vv124: OR2 port map(Z0 => v174, A0 => v175, A1 => K7);

    vv125: NAND2 port map(ZN0 => v107, A0 => v103, A1 => v104);
    vv126: NAND2 port map(ZN0 => v117, A0 => v113, A1 => v114);
    vv127: NAND2 port map(ZN0 => v127, A0 => v123, A1 => v124);
    vv128: NAND2 port map(ZN0 => v137, A0 => v133, A1 => v134);
    vv129: NAND2 port map(ZN0 => v147, A0 => v143, A1 => v144);
    vv130: NAND2 port map(ZN0 => v157, A0 => v153, A1 => v154);
    vv131: NAND2 port map(ZN0 => v167, A0 => v163, A1 => v164);
    vv132: NAND2 port map(ZN0 => v177, A0 => v173, A1 => v174);

    vv133: INV port map(ZN0 => v105, A0 => v106);
    vv134: INV port map(ZN0 => v115, A0 => v116);
    vv135: INV port map(ZN0 => v125, A0 => v126);
    vv136: INV port map(ZN0 => v135, A0 => v136);
    vv137: INV port map(ZN0 => v145, A0 => v146);
    vv138: INV port map(ZN0 => v155, A0 => v156);
    vv139: INV port map(ZN0 => v165, A0 => v166);
    vv140: INV port map(ZN0 => v175, A0 => v176);

    vv141: BUF port map(Z0 => Q0, A0 => v106);
    vv142: BUF port map(Z0 => Q1, A0 => v116);
    vv143: BUF port map(Z0 => Q2, A0 => v126);
    vv144: BUF port map(Z0 => Q3, A0 => v136);
    vv145: BUF port map(Z0 => Q4, A0 => v146);
    vv146: BUF port map(Z0 => Q5, A0 => v156);
    vv147: BUF port map(Z0 => Q6, A0 => v166);
    vv148: BUF port map(Z0 => Q7, A0 => v176);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK71 is
    port(Q0: OUT std_logic;
         J0: IN std_logic;
         K0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end FJK71;

architecture LATTICE_ARCH of FJK71 is
    signal v104: std_logic;
    signal v102: std_logic;
    signal v100: std_logic;
    signal v103: std_logic;
    signal v101: std_logic;
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
begin
    v111: FDE1
        port map(Q0 => v103,
                 D0 => v104,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v112: NAND2
        port map(ZN0 => v100,
                 A0 => v102,
                 A1 => J0);
    
    v113: OR2
        port map(Z0 => v101,
                 A0 => v102,
                 A1 => K0);
    
    v114: NAND2
        port map(ZN0 => v104,
                 A0 => v100,
                 A1 => v101);
    
    v115: INV
        port map(ZN0 => v102,
                 A0 => v103);
    
    v116: BUF
        port map(Z0 => Q0,
                 A0 => v103);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK71E is
    port(Q0: OUT std_logic;
         J0: IN std_logic;
         K0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end FJK71E;

architecture LATTICE_ARCH of FJK71E is
    signal v108: std_logic;
    signal v106: std_logic;
    signal v104: std_logic;
    signal v107: std_logic;
    signal v105: std_logic;
    
    component FDE1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : FDE1E use entity LAT_VHD.FDE1E(LATTICE_ARCH);
    
    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);
    
    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
begin
    v115: FDE1E
        port map(Q0 => v107,
                 D0 => v108,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    v116: NAND2
        port map(ZN0 => v104,
                 A0 => v106,
                 A1 => J0);
    
    v117: OR2
        port map(Z0 => v105,
                 A0 => v106,
                 A1 => K0);
    
    v118: NAND2
        port map(ZN0 => v108,
                 A0 => v104,
                 A1 => v105);
    
    v119: INV
        port map(ZN0 => v106,
                 A0 => v107);
    
    v120: BUF
        port map(Z0 => Q0,
                 A0 => v107);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK74 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         J0: IN std_logic;
         J1: IN std_logic;
         J2: IN std_logic;
         J3: IN std_logic;
         K0: IN std_logic;
         K1: IN std_logic;
         K2: IN std_logic;
         K3: IN std_logic;
         CLK: IN std_logic);
end FJK74;

architecture LATTICE_ARCH of FJK74 is
    signal v100,v101,v102,v103,v104 : std_logic;
    signal v110,v111,v112,v113,v114 : std_logic;
    signal v120,v121,v122,v123,v124 : std_logic;
    signal v130,v131,v132,v133,v134 : std_logic;

    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);

    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);

    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

begin
    vv100: FDE1 port map(Q0 => v103, D0 => v104, CLK => CLK, SD => SD, CD => CD);
    vv101: FDE1 port map(Q0 => v113, D0 => v114, CLK => CLK, SD => SD, CD => CD);
    vv102: FDE1 port map(Q0 => v123, D0 => v124, CLK => CLK, SD => SD, CD => CD);
    vv103: FDE1 port map(Q0 => v133, D0 => v134, CLK => CLK, SD => SD, CD => CD);

    vv110: NAND2 port map(ZN0 => v100, A0 => v102, A1 => J0);
    vv111: NAND2 port map(ZN0 => v110, A0 => v112, A1 => J1);
    vv112: NAND2 port map(ZN0 => v120, A0 => v122, A1 => J2);
    vv113: NAND2 port map(ZN0 => v130, A0 => v132, A1 => J3);

    vv120: OR2 port map(Z0 => v101, A0 => v102, A1 => K0);
    vv121: OR2 port map(Z0 => v111, A0 => v112, A1 => K1);
    vv122: OR2 port map(Z0 => v121, A0 => v122, A1 => K2);
    vv123: OR2 port map(Z0 => v131, A0 => v132, A1 => K3);

    vv130: NAND2 port map(ZN0 => v104, A0 => v100, A1 => v101);
    vv131: NAND2 port map(ZN0 => v114, A0 => v110, A1 => v111);
    vv132: NAND2 port map(ZN0 => v124, A0 => v120, A1 => v121);
    vv133: NAND2 port map(ZN0 => v134, A0 => v130, A1 => v131);

    vv140: INV port map(ZN0 => v102, A0 => v103);
    vv141: INV port map(ZN0 => v112, A0 => v113);
    vv142: INV port map(ZN0 => v122, A0 => v123);
    vv143: INV port map(ZN0 => v132, A0 => v133);

    vv150: BUF port map(Z0 => Q0, A0 => v103);
    vv151: BUF port map(Z0 => Q1, A0 => v113);
    vv152: BUF port map(Z0 => Q2, A0 => v123);
    vv153: BUF port map(Z0 => Q3, A0 => v133);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK74E is
    port(CD: IN std_logic;
	 SD: IN std_logic;
	 Q0: OUT std_logic;
	 Q1: OUT std_logic;
	 Q2: OUT std_logic;
	 Q3: OUT std_logic;
	 J0: IN std_logic;
	 J1: IN std_logic;
	 J2: IN std_logic;
	 J3: IN std_logic;
	 K0: IN std_logic;
	 K1: IN std_logic;
	 K2: IN std_logic;
	 K3: IN std_logic;
	 CLK: IN std_logic;
	 EN: IN std_logic);
end FJK74E;

architecture LATTICE_ARCH of FJK74E is
    signal v100,v101,v102,v103,v104 : std_logic;
    signal v110,v111,v112,v113,v114 : std_logic;
    signal v120,v121,v122,v123,v124 : std_logic;
    signal v130,v131,v132,v133,v134 : std_logic;

    component FDE1E
	port(Q0: OUT std_logic;
	     D0: IN std_logic;
	     CLK: IN std_logic;
	     SD: IN std_logic;
	     CD: IN std_logic;
	   EN: IN std_logic);
    end component;
    for all : FDE1E use entity LAT_VHD.FDE1E(LATTICE_ARCH);

    component NAND2
	port(ZN0: OUT std_logic;
	     A0: IN std_logic;
	     A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);

    component OR2
	port(Z0: OUT std_logic;
	     A0: IN std_logic;
	     A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);

    component INV
	port(ZN0: OUT std_logic;
	     A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
	port(Z0: OUT std_logic;
	     A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

begin
    vv100: FDE1E port map(Q0 => v103, D0 => v104, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv101: FDE1E port map(Q0 => v113, D0 => v114, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv102: FDE1E port map(Q0 => v123, D0 => v124, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv103: FDE1E port map(Q0 => v133, D0 => v134, CLK => CLK, SD => SD, CD => CD, EN => EN);

    vv110: NAND2 port map(ZN0 => v100, A0 => v102, A1 => J0);
    vv111: NAND2 port map(ZN0 => v110, A0 => v112, A1 => J1);
    vv112: NAND2 port map(ZN0 => v120, A0 => v122, A1 => J2);
    vv113: NAND2 port map(ZN0 => v130, A0 => v132, A1 => J3);

    vv120: OR2 port map(Z0 => v101, A0 => v102, A1 => K0);
    vv121: OR2 port map(Z0 => v111, A0 => v112, A1 => K1);
    vv122: OR2 port map(Z0 => v121, A0 => v122, A1 => K2);
    vv123: OR2 port map(Z0 => v131, A0 => v132, A1 => K3);

    vv130: NAND2 port map(ZN0 => v104, A0 => v100, A1 => v101);
    vv131: NAND2 port map(ZN0 => v114, A0 => v110, A1 => v111);
    vv132: NAND2 port map(ZN0 => v124, A0 => v120, A1 => v121);
    vv133: NAND2 port map(ZN0 => v134, A0 => v130, A1 => v131);

    vv140: INV port map(ZN0 => v102, A0 => v103);
    vv141: INV port map(ZN0 => v112, A0 => v113);
    vv142: INV port map(ZN0 => v122, A0 => v123);
    vv143: INV port map(ZN0 => v132, A0 => v133);

    vv150: BUF port map(Z0 => Q0, A0 => v103);
    vv151: BUF port map(Z0 => Q1, A0 => v113);
    vv152: BUF port map(Z0 => Q2, A0 => v123);
    vv153: BUF port map(Z0 => Q3, A0 => v133);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK78 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         J0: IN std_logic;
         J1: IN std_logic;
         J2: IN std_logic;
         J3: IN std_logic;
         J4: IN std_logic;
         J5: IN std_logic;
         J6: IN std_logic;
         J7: IN std_logic;
         K0: IN std_logic;
         K1: IN std_logic;
         K2: IN std_logic;
         K3: IN std_logic;
         K4: IN std_logic;
         K5: IN std_logic;
         K6: IN std_logic;
         K7: IN std_logic;
         CLK: IN std_logic);
end FJK78;

architecture LATTICE_ARCH of FJK78 is
    signal v100,v101,v102,v103,v104 : std_logic;
    signal v110,v111,v112,v113,v114 : std_logic;
    signal v120,v121,v122,v123,v124 : std_logic;
    signal v130,v131,v132,v133,v134 : std_logic;
    signal v140,v141,v142,v143,v144 : std_logic;
    signal v150,v151,v152,v153,v154 : std_logic;
    signal v160,v161,v162,v163,v164 : std_logic;
    signal v170,v171,v172,v173,v174 : std_logic;

    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);

    component NAND2
        port(ZN0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);

    component OR2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

begin
    vv100: FDE1 port map(Q0 => v103, D0 => v104, CLK => CLK, SD => SD, CD => CD);
    vv101: FDE1 port map(Q0 => v113, D0 => v114, CLK => CLK, SD => SD, CD => CD);
    vv102: FDE1 port map(Q0 => v123, D0 => v124, CLK => CLK, SD => SD, CD => CD);
    vv103: FDE1 port map(Q0 => v133, D0 => v134, CLK => CLK, SD => SD, CD => CD);
    vv104: FDE1 port map(Q0 => v143, D0 => v144, CLK => CLK, SD => SD, CD => CD);
    vv105: FDE1 port map(Q0 => v153, D0 => v154, CLK => CLK, SD => SD, CD => CD);
    vv106: FDE1 port map(Q0 => v163, D0 => v164, CLK => CLK, SD => SD, CD => CD);
    vv107: FDE1 port map(Q0 => v173, D0 => v174, CLK => CLK, SD => SD, CD => CD);

    vv110: NAND2 port map(ZN0 => v100, A0 => v102, A1 => J0);
    vv111: NAND2 port map(ZN0 => v110, A0 => v112, A1 => J1);
    vv112: NAND2 port map(ZN0 => v120, A0 => v122, A1 => J2);
    vv113: NAND2 port map(ZN0 => v130, A0 => v132, A1 => J3);
    vv114: NAND2 port map(ZN0 => v140, A0 => v142, A1 => J4);
    vv115: NAND2 port map(ZN0 => v150, A0 => v152, A1 => J5);
    vv116: NAND2 port map(ZN0 => v160, A0 => v162, A1 => J6);
    vv117: NAND2 port map(ZN0 => v170, A0 => v172, A1 => J7);

    vv120: OR2 port map(Z0 => v101, A0 => v102, A1 => K0);
    vv121: OR2 port map(Z0 => v111, A0 => v112, A1 => K1);
    vv122: OR2 port map(Z0 => v121, A0 => v122, A1 => K2);
    vv123: OR2 port map(Z0 => v131, A0 => v132, A1 => K3);
    vv124: OR2 port map(Z0 => v141, A0 => v142, A1 => K4);
    vv125: OR2 port map(Z0 => v151, A0 => v152, A1 => K5);
    vv126: OR2 port map(Z0 => v161, A0 => v162, A1 => K6);
    vv127: OR2 port map(Z0 => v171, A0 => v172, A1 => K7);

    vv130: NAND2 port map(ZN0 => v104, A0 => v100, A1 => v101);
    vv131: NAND2 port map(ZN0 => v114, A0 => v110, A1 => v111);
    vv132: NAND2 port map(ZN0 => v124, A0 => v120, A1 => v121);
    vv133: NAND2 port map(ZN0 => v134, A0 => v130, A1 => v131);
    vv134: NAND2 port map(ZN0 => v144, A0 => v140, A1 => v141);
    vv135: NAND2 port map(ZN0 => v154, A0 => v150, A1 => v151);
    vv136: NAND2 port map(ZN0 => v164, A0 => v160, A1 => v161);
    vv137: NAND2 port map(ZN0 => v174, A0 => v170, A1 => v171);

    vv140: INV port map(ZN0 => v102, A0 => v103);
    vv141: INV port map(ZN0 => v112, A0 => v113);
    vv142: INV port map(ZN0 => v122, A0 => v123);
    vv143: INV port map(ZN0 => v132, A0 => v133);
    vv144: INV port map(ZN0 => v142, A0 => v143);
    vv145: INV port map(ZN0 => v152, A0 => v153);
    vv146: INV port map(ZN0 => v162, A0 => v163);
    vv147: INV port map(ZN0 => v172, A0 => v173);

    vv150: BUF port map(Z0 => Q0, A0 => v103);
    vv151: BUF port map(Z0 => Q1, A0 => v113);
    vv152: BUF port map(Z0 => Q2, A0 => v123);
    vv153: BUF port map(Z0 => Q3, A0 => v133);
    vv154: BUF port map(Z0 => Q4, A0 => v143);
    vv155: BUF port map(Z0 => Q5, A0 => v153);
    vv156: BUF port map(Z0 => Q6, A0 => v163);
    vv157: BUF port map(Z0 => Q7, A0 => v173);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity FJK78 is
    port(CD: IN std_logic;
	 SD: IN std_logic;
	 Q0: OUT std_logic;
	 Q1: OUT std_logic;
	 Q2: OUT std_logic;
	 Q3: OUT std_logic;
	 Q4: OUT std_logic;
	 Q5: OUT std_logic;
	 Q6: OUT std_logic;
	 Q7: OUT std_logic;
	 J0: IN std_logic;
	 J1: IN std_logic;
	 J2: IN std_logic;
	 J3: IN std_logic;
	 J4: IN std_logic;
	 J5: IN std_logic;
	 J6: IN std_logic;
	 J7: IN std_logic;
	 K0: IN std_logic;
	 K1: IN std_logic;
	 K2: IN std_logic;
	 K3: IN std_logic;
	 K4: IN std_logic;
	 K5: IN std_logic;
	 K6: IN std_logic;
	 K7: IN std_logic;
	 CLK: IN std_logic;
	 EN: IN std_logic);
end FJK78;

architecture LATTICE_ARCH of FJK78 is
    signal v100,v101,v102,v103,v104 : std_logic;
    signal v110,v111,v112,v113,v114 : std_logic;
    signal v120,v121,v122,v123,v124 : std_logic;
    signal v130,v131,v132,v133,v134 : std_logic;
    signal v140,v141,v142,v143,v144 : std_logic;
    signal v150,v151,v152,v153,v154 : std_logic;
    signal v160,v161,v162,v163,v164 : std_logic;
    signal v170,v171,v172,v173,v174 : std_logic;

    component FDE1E
	port(Q0: OUT std_logic;
	     D0: IN std_logic;
	     CLK: IN std_logic;
	     SD: IN std_logic;
	     CD: IN std_logic;
	   EN: IN std_logic);
    end component;
    for all : FDE1E use entity LAT_VHD.FDE1E(LATTICE_ARCH);

    component NAND2
	port(ZN0: OUT std_logic;
	     A0: IN std_logic;
	     A1: IN std_logic);
    end component;
    for all : NAND2 use entity LAT_VHD.NAND2(LATTICE_ARCH);

    component OR2
	port(Z0: OUT std_logic;
	     A0: IN std_logic;
	     A1: IN std_logic);
    end component;
    for all : OR2 use entity LAT_VHD.OR2(LATTICE_ARCH);

    component INV
	port(ZN0: OUT std_logic;
	     A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
	port(Z0: OUT std_logic;
	     A0: IN std_logic);
    end component;
    for all : BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

begin
    vv100: FDE1E port map(Q0 => v103, D0 => v104, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv101: FDE1E port map(Q0 => v113, D0 => v114, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv102: FDE1E port map(Q0 => v123, D0 => v124, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv103: FDE1E port map(Q0 => v133, D0 => v134, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv104: FDE1E port map(Q0 => v143, D0 => v144, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv105: FDE1E port map(Q0 => v153, D0 => v154, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv106: FDE1E port map(Q0 => v163, D0 => v164, CLK => CLK, SD => SD, CD => CD, EN => EN);
    vv107: FDE1E port map(Q0 => v173, D0 => v174, CLK => CLK, SD => SD, CD => CD, EN => EN);

    vv110: NAND2 port map(ZN0 => v100, A0 => v102, A1 => J0);
    vv111: NAND2 port map(ZN0 => v110, A0 => v112, A1 => J1);
    vv112: NAND2 port map(ZN0 => v120, A0 => v122, A1 => J2);
    vv113: NAND2 port map(ZN0 => v130, A0 => v132, A1 => J3);
    vv114: NAND2 port map(ZN0 => v140, A0 => v142, A1 => J4);
    vv115: NAND2 port map(ZN0 => v150, A0 => v152, A1 => J5);
    vv116: NAND2 port map(ZN0 => v160, A0 => v162, A1 => J6);
    vv117: NAND2 port map(ZN0 => v170, A0 => v172, A1 => J7);

    vv120: OR2 port map(Z0 => v101, A0 => v102, A1 => K0);
    vv121: OR2 port map(Z0 => v111, A0 => v112, A1 => K1);
    vv122: OR2 port map(Z0 => v121, A0 => v122, A1 => K2);
    vv123: OR2 port map(Z0 => v131, A0 => v132, A1 => K3);
    vv124: OR2 port map(Z0 => v141, A0 => v142, A1 => K4);
    vv125: OR2 port map(Z0 => v151, A0 => v152, A1 => K5);
    vv126: OR2 port map(Z0 => v161, A0 => v162, A1 => K6);
    vv127: OR2 port map(Z0 => v171, A0 => v172, A1 => K7);

    vv130: NAND2 port map(ZN0 => v104, A0 => v100, A1 => v101);
    vv131: NAND2 port map(ZN0 => v114, A0 => v110, A1 => v111);
    vv132: NAND2 port map(ZN0 => v124, A0 => v120, A1 => v121);
    vv133: NAND2 port map(ZN0 => v134, A0 => v130, A1 => v131);
    vv134: NAND2 port map(ZN0 => v144, A0 => v140, A1 => v141);
    vv135: NAND2 port map(ZN0 => v154, A0 => v150, A1 => v151);
    vv136: NAND2 port map(ZN0 => v164, A0 => v160, A1 => v161);
    vv137: NAND2 port map(ZN0 => v174, A0 => v170, A1 => v171);

    vv140: INV port map(ZN0 => v102, A0 => v103);
    vv141: INV port map(ZN0 => v112, A0 => v113);
    vv142: INV port map(ZN0 => v122, A0 => v123);
    vv143: INV port map(ZN0 => v132, A0 => v133);
    vv144: INV port map(ZN0 => v142, A0 => v143);
    vv145: INV port map(ZN0 => v152, A0 => v153);
    vv146: INV port map(ZN0 => v162, A0 => v163);
    vv147: INV port map(ZN0 => v172, A0 => v173);

    vv150: BUF port map(Z0 => Q0, A0 => v103);
    vv151: BUF port map(Z0 => Q1, A0 => v113);
    vv152: BUF port map(Z0 => Q2, A0 => v123);
    vv153: BUF port map(Z0 => Q3, A0 => v133);
    vv154: BUF port map(Z0 => Q4, A0 => v143);
    vv155: BUF port map(Z0 => Q5, A0 => v153);
    vv156: BUF port map(Z0 => Q6, A0 => v163);
    vv157: BUF port map(Z0 => Q7, A0 => v173);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID11E is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic);
end ID11E;

architecture LATTICE_ARCH of ID11E is
    signal v106: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);
    
begin
    v109: XINPUT
        port map(Z0 => v106,
                 XI0 => XI0);
    
    v110: XDFF1E
        port map(Q0 => Q0,
                 D0 => v106,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID14E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic);
end ID14E;

architecture LATTICE_ARCH of ID14E is
    signal v106, v116, v126, v136: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);

    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);

begin

    v100: XINPUT port map(Z0 => v106, XI0 => XI0);
    v101: XINPUT port map(Z0 => v116, XI0 => XI1);
    v102: XINPUT port map(Z0 => v126, XI0 => XI2);
    v103: XINPUT port map(Z0 => v136, XI0 => XI3);

    v110: XDFF1E port map(Q0 => Q0, D0 => v106, CLK => CLK, EN => EN);
    v111: XDFF1E port map(Q0 => Q1, D0 => v116, CLK => CLK, EN => EN);
    v112: XDFF1E port map(Q0 => Q2, D0 => v126, CLK => CLK, EN => EN);
    v113: XDFF1E port map(Q0 => Q3, D0 => v136, CLK => CLK, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID31 is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic);
end ID31;

architecture LATTICE_ARCH of ID31 is
    signal v103: std_logic;
    
    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
begin
    v106: XDFF2
        port map(Q0 => Q0,
                 D0 => v103,
                 CLK => CLK,
                 CD => CD);
    
    v107: XINPUT
        port map(Z0 => v103,
                 XI0 => XI0);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID31E is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic);
end ID31E;

architecture LATTICE_ARCH of ID31E is
    signal v107: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);
    
begin
    v110: XINPUT
        port map(Z0 => v107,
                 XI0 => XI0);
    
    v111: XDFF2E
        port map(Q0 => Q0,
                 D0 => v107,
                 CLK => CLK,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID34 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic);
end ID34;

architecture LATTICE_ARCH of ID34 is
    signal v103, v113, v123, v133: std_logic;

    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);

begin

    vv100: XDFF2 port map(Q0 => Q0, D0 => v103, CLK => CLK, CD => CD);
    vv101: XDFF2 port map(Q0 => Q1, D0 => v113, CLK => CLK, CD => CD);
    vv102: XDFF2 port map(Q0 => Q2, D0 => v123, CLK => CLK, CD => CD);
    vv103: XDFF2 port map(Q0 => Q3, D0 => v133, CLK => CLK, CD => CD);

    vv110: XINPUT port map(Z0 => v103, XI0 => XI0);
    vv111: XINPUT port map(Z0 => v113, XI0 => XI1);
    vv112: XINPUT port map(Z0 => v123, XI0 => XI2);
    vv113: XINPUT port map(Z0 => v133, XI0 => XI3);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID34E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic);
end ID34E;

architecture LATTICE_ARCH of ID34E is
    signal v107, v117, v127, v137: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
        end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
  
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);

begin

    v100: XINPUT port map(Z0 => v107, XI0 => XI0);
    v101: XINPUT port map(Z0 => v117, XI0 => XI1);
    v102: XINPUT port map(Z0 => v127, XI0 => XI2);
    v103: XINPUT port map(Z0 => v137, XI0 => XI3);

    v110: XDFF2E port map(Q0 => Q0, D0 => v107, CLK => CLK, CD => CD, EN => EN);
    v111: XDFF2E port map(Q0 => Q1, D0 => v117, CLK => CLK, CD => CD, EN => EN);
    v112: XDFF2E port map(Q0 => Q2, D0 => v127, CLK => CLK, CD => CD, EN => EN);
    v113: XDFF2E port map(Q0 => Q3, D0 => v137, CLK => CLK, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID41 is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic);
end ID41;

architecture LATTICE_ARCH of ID41 is
    signal v103: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);
    
begin
    v106: XINPUT
        port map(Z0 => v103,
                 XI0 => XI0);
    
    v107: XDFF3
        port map(Q0 => Q0,
                 D0 => v103,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID41E is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end ID41E;

architecture LATTICE_ARCH of ID41E is
    signal v107: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);
    
begin
    v110: XINPUT
        port map(Z0 => v107,
                 XI0 => XI0);
    
    v111: XDFF3E
        port map(Q0 => Q0,
                 D0 => v107,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID44 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic);
end ID44;

architecture LATTICE_ARCH of ID44 is
    signal v103, v113, v123, v133: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);

    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);

begin

    vv100: XINPUT port map(Z0 => v103, XI0 => XI0);
    vv101: XINPUT port map(Z0 => v113, XI0 => XI1);
    vv102: XINPUT port map(Z0 => v123, XI0 => XI2);
    vv103: XINPUT port map(Z0 => v133, XI0 => XI3);

    vv110: XDFF3 port map(Q0 => Q0, D0 => v103, CLK => CLK, SD => SD);
    vv111: XDFF3 port map(Q0 => Q1, D0 => v113, CLK => CLK, SD => SD);
    vv112: XDFF3 port map(Q0 => Q2, D0 => v123, CLK => CLK, SD => SD);
    vv113: XDFF3 port map(Q0 => Q3, D0 => v133, CLK => CLK, SD => SD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID44E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end ID44E;

architecture LATTICE_ARCH of ID44E is
    signal v107, v117, v127, v137: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
   
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);

begin

    v100: XINPUT port map(Z0 => v107, XI0 => XI0);
    v101: XINPUT port map(Z0 => v117, XI0 => XI1);
    v102: XINPUT port map(Z0 => v127, XI0 => XI2);
    v103: XINPUT port map(Z0 => v137, XI0 => XI3);

    v110: XDFF3E port map(Q0 => Q0, D0 => v107, CLK => CLK, SD => SD, EN => EN);
    v111: XDFF3E port map(Q0 => Q1, D0 => v117, CLK => CLK, SD => SD, EN => EN);
    v112: XDFF3E port map(Q0 => Q2, D0 => v127, CLK => CLK, SD => SD, EN => EN);
    v113: XDFF3E port map(Q0 => Q3, D0 => v137, CLK => CLK, SD => SD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID51 is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end ID51;

architecture LATTICE_ARCH of ID51 is
    signal v100: std_logic;
    
    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
begin
    v103: XDFF4
        port map(Q0 => Q0,
                 D0 => v100,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v104: XINPUT
        port map(Z0 => v100,
                 XI0 => XI0);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID51E is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end ID51E;

architecture LATTICE_ARCH of ID51E is
    signal v104: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);
    
begin
    v107: XINPUT
        port map(Z0 => v104,
                 XI0 => XI0);
    
    v108: XDFF4E
        port map(Q0 => Q0,
                 D0 => v104,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID54 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end ID54;

architecture LATTICE_ARCH of ID54 is
    signal v100, v110, v120, v130: std_logic;

    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
   
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);

begin

    vv100: XDFF4 port map(Q0 => Q0, D0 => v100, CLK => CLK, SD => SD, CD => CD);
    vv101: XDFF4 port map(Q0 => Q1, D0 => v110, CLK => CLK, SD => SD, CD => CD);
    vv102: XDFF4 port map(Q0 => Q2, D0 => v120, CLK => CLK, SD => SD, CD => CD);
    vv103: XDFF4 port map(Q0 => Q3, D0 => v130, CLK => CLK, SD => SD, CD => CD);

    vv110: XINPUT port map(Z0 => v100, XI0 => XI0);
    vv111: XINPUT port map(Z0 => v110, XI0 => XI1);
    vv112: XINPUT port map(Z0 => v120, XI0 => XI2);
    vv113: XINPUT port map(Z0 => v130, XI0 => XI3);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ID54E is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end ID54E;

architecture LATTICE_ARCH of ID54E is
    signal v104, v114, v124, v134: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
   
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);

begin

    v100: XINPUT port map(Z0 => v104, XI0 => XI0);
    v101: XINPUT port map(Z0 => v114, XI0 => XI1);
    v102: XINPUT port map(Z0 => v124, XI0 => XI2);
    v103: XINPUT port map(Z0 => v134, XI0 => XI3);

    v110: XDFF4E port map(Q0 => Q0, D0 => v104, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v111: XDFF4E port map(Q0 => Q1, D0 => v114, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v112: XDFF4E port map(Q0 => Q2, D0 => v124, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v113: XDFF4E port map(Q0 => Q3, D0 => v134, CLK => CLK, SD => SD, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IL31 is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic);
end IL31;

architecture LATTICE_ARCH of IL31 is
    signal v103: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);
    
begin
    v106: XINPUT
        port map(Z0 => v103,
                 XI0 => XI0);
    
    v107: XDL2
        port map(Q0 => Q0,
                 D0 => v103,
                 G => G,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IL34 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic);
end IL34;

architecture LATTICE_ARCH of IL34 is
    signal v103, v113, v123, v133: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);

    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);

begin

    vv100: XINPUT port map(Z0 => v103, XI0 => XI0);
    vv101: XINPUT port map(Z0 => v113, XI0 => XI1);
    vv102: XINPUT port map(Z0 => v123, XI0 => XI2);
    vv103: XINPUT port map(Z0 => v133, XI0 => XI3);

    vv110: XDL2 port map(Q0 => Q0, D0 => v103, G => G, CD => CD);
    vv111: XDL2 port map(Q0 => Q1, D0 => v113, G => G, CD => CD);
    vv112: XDL2 port map(Q0 => Q2, D0 => v123, G => G, CD => CD);
    vv113: XDL2 port map(Q0 => Q3, D0 => v133, G => G, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IL41 is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic);
end IL41;

architecture LATTICE_ARCH of IL41 is
    signal v103: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);
    
begin
    v106: XINPUT
        port map(Z0 => v103,
                 XI0 => XI0);
    
    v107: XDL3
        port map(Q0 => Q0,
                 D0 => v103,
                 G => G,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IL44 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic);
end IL44;

architecture LATTICE_ARCH of IL44 is
    signal v103, v113, v123, v133: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);

    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);

begin

    vv100: XINPUT port map(Z0 => v103, XI0 => XI0);
    vv101: XINPUT port map(Z0 => v113, XI0 => XI1);
    vv102: XINPUT port map(Z0 => v123, XI0 => XI2);
    vv103: XINPUT port map(Z0 => v133, XI0 => XI3);

    vv110: XDL3 port map(Q0 => Q0, D0 => v103, G => G, SD => SD);
    vv111: XDL3 port map(Q0 => Q1, D0 => v113, G => G, SD => SD);
    vv112: XDL3 port map(Q0 => Q2, D0 => v123, G => G, SD => SD);
    vv113: XDL3 port map(Q0 => Q3, D0 => v133, G => G, SD => SD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IL51 is
    port(Q0: OUT std_logic;
         XI0: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end IL51;

architecture LATTICE_ARCH of IL51 is
    signal v101: std_logic;
    
    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
    
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
    
begin
    v104: XINPUT
        port map(Z0 => v101,
                 XI0 => XI0);
    
    v105: XDL4
        port map(Q0 => Q0,
                 D0 => v101,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IL54 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         XI0: IN std_logic;
         XI1: IN std_logic;
         XI2: IN std_logic;
         XI3: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic;
         SD: IN std_logic);
end IL54;

architecture LATTICE_ARCH of IL54 is
    signal v101, v111, v121, v131: std_logic;

    component XINPUT
        port(Z0: OUT std_logic;
             XI0: IN std_logic);
    end component;
    for all : XINPUT use entity LAT_VHD.XINPUT(LATTICE_ARCH);
   
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);

begin

    vv100: XINPUT port map(Z0 => v101, XI0 => XI0);
    vv101: XINPUT port map(Z0 => v111, XI0 => XI1);
    vv102: XINPUT port map(Z0 => v121, XI0 => XI2);
    vv103: XINPUT port map(Z0 => v131, XI0 => XI3);

    vv110: XDL4 port map(Q0 => Q0, D0 => v101, G => G, SD => SD, CD => CD);
    vv111: XDL4 port map(Q0 => Q1, D0 => v111, G => G, SD => SD, CD => CD);
    vv112: XDL4 port map(Q0 => Q2, D0 => v121, G => G, SD => SD, CD => CD);
    vv113: XDL4 port map(Q0 => Q3, D0 => v131, G => G, SD => SD, CD => CD);

end LATTICE_ARCH;
Library IEEE;
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IT14 is
    port(OE: IN std_logic;
         O0: OUT std_logic;
         O1: OUT std_logic;
         O2: OUT std_logic;
         O3: OUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic);
end IT14;

architecture LATTICE_ARCH of IT14 is
    
    component IT11
        port(O0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);
    
begin
    v105: IT11
        port map(O0 => O0,
                 A0 => A0,
                 OE => OE);
    
    v106: IT11
        port map(O0 => O1,
                 A0 => A1,
                 OE => OE);
    
    v107: IT11
        port map(O0 => O2,
                 A0 => A2,
                 OE => OE);
    
    v108: IT11
        port map(O0 => O3,
                 A0 => A3,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IT18 is
    port(OE: IN std_logic;
         O0: OUT std_logic;
         O1: OUT std_logic;
         O2: OUT std_logic;
         O3: OUT std_logic;
         O4: OUT std_logic;
         O5: OUT std_logic;
         O6: OUT std_logic;
         O7: OUT std_logic;
         A0: IN std_logic;
         A1: IN std_logic;
         A2: IN std_logic;
         A3: IN std_logic;
         A4: IN std_logic;
         A5: IN std_logic;
         A6: IN std_logic;
         A7: IN std_logic);
end IT18;

architecture LATTICE_ARCH of IT18 is
    
    component IT11
        port(O0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);
    
begin
    v109: IT11
        port map(O0 => O0,
                 A0 => A0,
                 OE => OE);
    
    v110: IT11
        port map(O0 => O1,
                 A0 => A1,
                 OE => OE);
    
    v111: IT11
        port map(O0 => O2,
                 A0 => A2,
                 OE => OE);
    
    v112: IT11
        port map(O0 => O3,
                 A0 => A3,
                 OE => OE);
    
    v113: IT11
        port map(O0 => O4,
                 A0 => A4,
                 OE => OE);
    
    v114: IT11
        port map(O0 => O6,
                 A0 => A6,
                 OE => OE);
    
    v115: IT11
        port map(O0 => O7,
                 A0 => A7,
                 OE => OE);
    
    v116: IT11
        port map(O0 => O5,
                 A0 => A5,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IT21 is
    port(O0: OUT std_logic;
         A0: IN std_logic;
         OE: IN std_logic);
end IT21;

architecture LATTICE_ARCH of IT21 is
    signal v101: std_logic;
    
    component IT11
        port(O0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
begin
    v104: IT11
        port map(O0 => O0,
                 A0 => A0,
                 OE => v101);
    
    v105: INV
        port map(ZN0 => v101,
                 A0 => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IT24 is
    port(OE: IN std_logic;
	 O0: OUT std_logic;
	 O1: OUT std_logic;
	 O2: OUT std_logic;
	 O3: OUT std_logic;
	 A0: IN std_logic;
	 A1: IN std_logic;
	 A2: IN std_logic;
	 A3: IN std_logic);
end IT24;

architecture LATTICE_ARCH of IT24 is
    signal v101 : std_logic;
    
    component IT11
	port(O0: OUT std_logic;
	     A0: IN std_logic;
	     OE: IN std_logic);
    end component;
    for all : IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);
    
    component INV
	port(ZN0: OUT std_logic;
	      A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);

begin
    v106: IT11
	port map(O0 => O0,
		 A0 => A0,
		 OE => v101);
    
    v107: IT11
	port map(O0 => O1,
		 A0 => A1,
		 OE => v101);
    
    v108: IT11
	port map(O0 => O2,
		 A0 => A2,
		 OE => v101);
    
    v109: IT11
	port map(O0 => O3,
		 A0 => A3,
		 OE => v101);
    
    v110: INV
	port map(ZN0 => v101,
		  A0 => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity IT28 is
    port(OE: IN std_logic;
	 O0: OUT std_logic;
	 O1: OUT std_logic;
	 O2: OUT std_logic;
	 O3: OUT std_logic;
	 O4: OUT std_logic;
	 O5: OUT std_logic;
	 O6: OUT std_logic;
	 O7: OUT std_logic;
	 A0: IN std_logic;
	 A1: IN std_logic;
	 A2: IN std_logic;
	 A3: IN std_logic;
	 A4: IN std_logic;
	 A5: IN std_logic;
	 A6: IN std_logic;
	 A7: IN std_logic);
end IT28;

architecture LATTICE_ARCH of IT28 is
    signal v101 : std_logic;
    
    component IT11
	port(O0: OUT std_logic;
	     A0: IN std_logic;
	     OE: IN std_logic);
    end component;
    for all : IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);

    component INV
	port(ZN0: OUT std_logic;
	      A0: IN std_logic);
    end component;
    for all : INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
begin
    v110: IT11
	port map(O0 => O0,
		 A0 => A0,
		 OE => v101);
    
    v111: IT11
	port map(O0 => O1,
		 A0 => A1,
		 OE => v101);
    
    v112: IT11
	port map(O0 => O2,
		 A0 => A2,
		 OE => v101);
    
    v113: IT11
	port map(O0 => O3,
		 A0 => A3,
		 OE => v101);
    
    v114: IT11
	port map(O0 => O4,
		 A0 => A4,
		 OE => v101);
    
    v115: IT11
	port map(O0 => O5,
		 A0 => A5,
		 OE => v101);
    
    v116: IT11
	port map(O0 => O6,
		 A0 => A6,
		 OE => v101);
    
    v117: IT11
	port map(O0 => O7,
		 A0 => A7,
		 OE => v101);
    
    v118: INV
	port map(ZN0 => v101,
		  A0 => OE);
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI14 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic);
end LDI14;

architecture LATTICE_ARCH of LDI14 is
    
    component LDI11
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: LDI11 use entity LAT_VHD.LDI11(LATTICE_ARCH);
    
begin
    v106: LDI11
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G);
    
    v107: LDI11
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G);
    
    v108: LDI11
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G);
    
    v109: LDI11
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI18 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         G: IN std_logic);
end LDI18;

architecture LATTICE_ARCH of LDI18 is
    
    component LDI11
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: LDI11 use entity LAT_VHD.LDI11(LATTICE_ARCH);
    
begin
    v110: LDI11
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G);
    
    v111: LDI11
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G);
    
    v112: LDI11
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G);
    
    v113: LDI11
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G);
    
    v114: LDI11
        port map(Q0 => Q4,
                 D0 => D4,
                 G => G);
    
    v115: LDI11
        port map(Q0 => Q5,
                 D0 => D5,
                 G => G);
    
    v116: LDI11
        port map(Q0 => Q6,
                 D0 => D6,
                 G => G);
    
    v117: LDI11
        port map(Q0 => Q7,
                 D0 => D7,
                 G => G);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI24 is
    port(CD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic);
end LDI24;

architecture LATTICE_ARCH of LDI24 is
    
    component LDI21
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: LDI21 use entity LAT_VHD.LDI21(LATTICE_ARCH);
    
begin
    v107: LDI21
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G,
                 CD => CD);
    
    v108: LDI21
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G,
                 CD => CD);
    
    v109: LDI21
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G,
                 CD => CD);
    
    v110: LDI21
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI28 is
    port(CD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         G: IN std_logic);
end LDI28;

architecture LATTICE_ARCH of LDI28 is
    
    component LDI21
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: LDI21 use entity LAT_VHD.LDI21(LATTICE_ARCH);
    
begin
    v111: LDI21
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G,
                 CD => CD);
    
    v112: LDI21
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G,
                 CD => CD);
    
    v113: LDI21
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G,
                 CD => CD);
    
    v114: LDI21
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G,
                 CD => CD);
    
    v115: LDI21
        port map(Q0 => Q4,
                 D0 => D4,
                 G => G,
                 CD => CD);
    
    v116: LDI21
        port map(Q0 => Q5,
                 D0 => D5,
                 G => G,
                 CD => CD);
    
    v117: LDI21
        port map(Q0 => Q6,
                 D0 => D6,
                 G => G,
                 CD => CD);
    
    v118: LDI21
        port map(Q0 => Q7,
                 D0 => D7,
                 G => G,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI34 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic);
end LDI34;

architecture LATTICE_ARCH of LDI34 is
    
    component LDI31
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: LDI31 use entity LAT_VHD.LDI31(LATTICE_ARCH);
    
begin
    v107: LDI31
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G,
                 SD => SD);
    
    v108: LDI31
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G,
                 SD => SD);
    
    v109: LDI31
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G,
                 SD => SD);
    
    v110: LDI31
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI38 is
    port(SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         G: IN std_logic);
end LDI38;

architecture LATTICE_ARCH of LDI38 is
    
    component LDI31
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: LDI31 use entity LAT_VHD.LDI31(LATTICE_ARCH);
    
begin
    v111: LDI31
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G,
                 SD => SD);
    
    v112: LDI31
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G,
                 SD => SD);
    
    v113: LDI31
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G,
                 SD => SD);
    
    v114: LDI31
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G,
                 SD => SD);
    
    v115: LDI31
        port map(Q0 => Q4,
                 D0 => D4,
                 G => G,
                 SD => SD);
    
    v116: LDI31
        port map(Q0 => Q5,
                 D0 => D5,
                 G => G,
                 SD => SD);
    
    v117: LDI31
        port map(Q0 => Q6,
                 D0 => D6,
                 G => G,
                 SD => SD);
    
    v118: LDI31
        port map(Q0 => Q7,
                 D0 => D7,
                 G => G,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI44 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic);
end LDI44;

architecture LATTICE_ARCH of LDI44 is
    
    component LDI41
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: LDI41 use entity LAT_VHD.LDI41(LATTICE_ARCH);
    
begin
    v104: LDI41
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v105: LDI41
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v106: LDI41
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v107: LDI41
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity LDI48 is
    port(CD: IN std_logic;
         SD: IN std_logic;
         Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         G: IN std_logic);
end LDI48;

architecture LATTICE_ARCH of LDI48 is
    
    component LDI41
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: LDI41 use entity LAT_VHD.LDI41(LATTICE_ARCH);
    
begin
    v108: LDI41
        port map(Q0 => Q0,
                 D0 => D0,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v109: LDI41
        port map(Q0 => Q1,
                 D0 => D1,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v110: LDI41
        port map(Q0 => Q2,
                 D0 => D2,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v111: LDI41
        port map(Q0 => Q3,
                 D0 => D3,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v112: LDI41
        port map(Q0 => Q4,
                 D0 => D4,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v113: LDI41
        port map(Q0 => Q5,
                 D0 => D5,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v114: LDI41
        port map(Q0 => Q6,
                 D0 => D6,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v115: LDI41
        port map(Q0 => Q7,
                 D0 => D7,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD11 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic);
end OD11;

architecture LATTICE_ARCH of OD11 is
    
    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);
    
begin
    v101: XDFF1
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD11E is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic);
end OD11E;

architecture LATTICE_ARCH of OD11E is
    
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);
    
begin
    v107: XDFF1E
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD14 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic);
end OD14;

architecture LATTICE_ARCH of OD14 is

    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);

begin
    v100: XDFF1 port map(Q0 => XQ0, D0 => D0, CLK => CLK);
    v101: XDFF1 port map(Q0 => XQ1, D0 => D1, CLK => CLK);
    v102: XDFF1 port map(Q0 => XQ2, D0 => D2, CLK => CLK);
    v103: XDFF1 port map(Q0 => XQ3, D0 => D3, CLK => CLK);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD14E is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic);
end OD14E;

architecture LATTICE_ARCH of OD14E is

    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);

begin
    v100: XDFF1E port map(Q0 => XQ0, D0 => D0, CLK => CLK, EN => EN);
    v101: XDFF1E port map(Q0 => XQ1, D0 => D1, CLK => CLK, EN => EN);
    v102: XDFF1E port map(Q0 => XQ2, D0 => D2, CLK => CLK, EN => EN);
    v103: XDFF1E port map(Q0 => XQ3, D0 => D3, CLK => CLK, EN => EN);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD21 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic);
end OD21;

architecture LATTICE_ARCH of OD21 is
    signal v100: std_logic;
    
    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
begin
    v103: XDFF1
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => v100);
    
    v104: INV
        port map(ZN0 => v100,
                 A0 => CLK);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD24 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic);
end OD24;

architecture LATTICE_ARCH of OD24 is
    signal v100: std_logic;

    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);

begin

    vv100: XDFF1 port map(Q0 => XQ0, D0 => D0, CLK => v100);
    vv101: XDFF1 port map(Q0 => XQ1, D0 => D1, CLK => v100);
    vv102: XDFF1 port map(Q0 => XQ2, D0 => D2, CLK => v100);
    vv103: XDFF1 port map(Q0 => XQ3, D0 => D3, CLK => v100);

    v110: INV port map(ZN0 => v100, A0 => CLK);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD31 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic);
end OD31;

architecture LATTICE_ARCH of OD31 is
    
    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);
    
begin
    v104: XDFF2
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD31E is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic);
end OD31E;

architecture LATTICE_ARCH of OD31E is
    
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);
    
begin
    v108: XDFF2E
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD34 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic);
end OD34;

architecture LATTICE_ARCH of OD34 is

    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);

begin
    v100: XDFF2 port map(Q0 => XQ0, D0 => D0, CLK => CLK, CD => CD);
    v101: XDFF2 port map(Q0 => XQ1, D0 => D1, CLK => CLK, CD => CD);
    v102: XDFF2 port map(Q0 => XQ2, D0 => D2, CLK => CLK, CD => CD);
    v103: XDFF2 port map(Q0 => XQ3, D0 => D3, CLK => CLK, CD => CD);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD34E is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic);
end OD34E;

architecture LATTICE_ARCH of OD34E is

    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);

begin
    v100: XDFF2E port map(Q0 => XQ0, D0 => D0, CLK => CLK, CD => CD, EN => EN);
    v101: XDFF2E port map(Q0 => XQ1, D0 => D1, CLK => CLK, CD => CD, EN => EN);
    v102: XDFF2E port map(Q0 => XQ2, D0 => D2, CLK => CLK, CD => CD, EN => EN);
    v103: XDFF2E port map(Q0 => XQ3, D0 => D3, CLK => CLK, CD => CD, EN => EN);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD41 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic);
end OD41;

architecture LATTICE_ARCH of OD41 is
    
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);
    
begin
    v104: XDFF3
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD41E is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end OD41E;

architecture LATTICE_ARCH of OD41E is
    
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);
    
begin
    v108: XDFF3E
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD44 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic);
end OD44;

architecture LATTICE_ARCH of OD44 is

    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);

begin
    v100: XDFF3 port map(Q0 => XQ0, D0 => D0, CLK => CLK, SD => SD);
    v101: XDFF3 port map(Q0 => XQ1, D0 => D1, CLK => CLK, SD => SD);
    v102: XDFF3 port map(Q0 => XQ2, D0 => D2, CLK => CLK, SD => SD);
    v103: XDFF3 port map(Q0 => XQ3, D0 => D3, CLK => CLK, SD => SD);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD44E is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic);
end OD44E;

architecture LATTICE_ARCH of OD44E is

    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);

begin
    v100: XDFF3E port map(Q0 => XQ0, D0 => D0, CLK => CLK, SD => SD, EN => EN);
    v101: XDFF3E port map(Q0 => XQ1, D0 => D1, CLK => CLK, SD => SD, EN => EN);
    v102: XDFF3E port map(Q0 => XQ2, D0 => D2, CLK => CLK, SD => SD, EN => EN);
    v103: XDFF3E port map(Q0 => XQ3, D0 => D3, CLK => CLK, SD => SD, EN => EN);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD51 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic);
end OD51;

architecture LATTICE_ARCH of OD51 is
    
    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
    
begin
    v101: XDFF4
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD51E is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic);
end OD51E;

architecture LATTICE_ARCH of OD51E is
    
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);
    
begin
    v105: XDFF4E
        port map(Q0 => XQ0,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD54 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic);
end OD54;

architecture LATTICE_ARCH of OD54 is

    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);

begin
    v100: XDFF4 port map(Q0 => XQ0, D0 => D0, CLK => CLK, SD => SD, CD => CD);
    v101: XDFF4 port map(Q0 => XQ1, D0 => D1, CLK => CLK, SD => SD, CD => CD);
    v102: XDFF4 port map(Q0 => XQ2, D0 => D2, CLK => CLK, SD => SD, CD => CD);
    v103: XDFF4 port map(Q0 => XQ3, D0 => D3, CLK => CLK, SD => SD, CD => CD);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OD54E is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic);
end OD54E;

architecture LATTICE_ARCH of OD54E is

    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all: XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);

begin
    v100: XDFF4E port map(Q0 => XQ0, D0 => D0, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v101: XDFF4E port map(Q0 => XQ1, D0 => D1, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v102: XDFF4E port map(Q0 => XQ2, D0 => D2, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v103: XDFF4E port map(Q0 => XQ3, D0 => D3, CLK => CLK, SD => SD, CD => CD, EN => EN);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT11 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end ODT11;

architecture LATTICE_ARCH of ODT11 is
    signal v101: std_logic;
    
    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v104: XDFF1
        port map(Q0 => v101,
                 D0 => D0,
                 CLK => CLK);
    
    v105: XTRI1
        port map(XO0 => XO0,
                 A0 => v101,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT11E is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end ODT11E;

architecture LATTICE_ARCH of ODT11E is
    signal v107: std_logic;
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);
    
begin
    v110: XTRI1
        port map(XO0 => XO0,
                 A0 => v107,
                 OE => OE);
    
    v111: XDFF1E
        port map(Q0 => v107,
                 D0 => D0,
                 CLK => CLK,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT14 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         OE: IN std_logic);
end ODT14;

architecture LATTICE_ARCH of ODT14 is
    signal v101, v111, v121, v131: std_logic;

    component XDFF1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic);
    end component;
    for all: XDFF1 use entity LAT_VHD.XDFF1(LATTICE_ARCH);

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    vv100: XDFF1 port map(Q0 => v101, D0 => D0, CLK => CLK);
    vv101: XDFF1 port map(Q0 => v111, D0 => D1, CLK => CLK);
    vv102: XDFF1 port map(Q0 => v121, D0 => D2, CLK => CLK);
    vv103: XDFF1 port map(Q0 => v131, D0 => D3, CLK => CLK);

    vv110: XTRI1 port map(XO0 => XO0, A0 => v101, OE => OE);
    vv111: XTRI1 port map(XO0 => XO1, A0 => v111, OE => OE);
    vv112: XTRI1 port map(XO0 => XO2, A0 => v121, OE => OE);
    vv113: XTRI1 port map(XO0 => XO3, A0 => v131, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT14E is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end ODT14E;

architecture LATTICE_ARCH of ODT14E is
    signal v107, v117, v127, v137: std_logic;
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
      
    component XDFF1E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF1E use entity LAT_VHD.XDFF1E(LATTICE_ARCH);

begin

    v100: XTRI1 port map(XO0 => XO0, A0 => v107, OE => OE);
    v101: XTRI1 port map(XO0 => XO1, A0 => v117, OE => OE);
    v102: XTRI1 port map(XO0 => XO2, A0 => v127, OE => OE);
    v103: XTRI1 port map(XO0 => XO3, A0 => v137, OE => OE);

    v110: XDFF1E port map(Q0 => v107, D0 => D0, CLK => CLK, EN => EN);
    v111: XDFF1E port map(Q0 => v117, D0 => D1, CLK => CLK, EN => EN);
    v112: XDFF1E port map(Q0 => v127, D0 => D2, CLK => CLK, EN => EN);
    v113: XDFF1E port map(Q0 => v137, D0 => D3, CLK => CLK, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT21 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT21;

architecture LATTICE_ARCH of ODT21 is
    signal v104: std_logic;
    
    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v107: XDFF2
        port map(Q0 => v104,
                 D0 => D0,
                 CLK => CLK,
                 CD => CD);
    
    v108: XTRI1
        port map(XO0 => XO0,
                 A0 => v104,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT21E is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT21E;

architecture LATTICE_ARCH of ODT21E is
    signal v108: std_logic;
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);
    
begin
    v111: XTRI1
        port map(XO0 => XO0,
                 A0 => v108,
                 OE => OE);
    
    v112: XDFF2E
        port map(Q0 => v108,
                 D0 => D0,
                 CLK => CLK,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT24 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT24;

architecture LATTICE_ARCH of ODT24 is
    signal v104, v114, v124, v134: std_logic;

    component XDFF2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF2 use entity LAT_VHD.XDFF2(LATTICE_ARCH);

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    vv101: XDFF2 port map(Q0 => v104, D0 => D0, CLK => CLK, CD => CD);
    vv102: XDFF2 port map(Q0 => v114, D0 => D1, CLK => CLK, CD => CD);
    vv103: XDFF2 port map(Q0 => v124, D0 => D2, CLK => CLK, CD => CD);
    vv104: XDFF2 port map(Q0 => v134, D0 => D3, CLK => CLK, CD => CD);

    vv111: XTRI1 port map(XO0 => XO0, A0 => v104, OE => OE);
    vv112: XTRI1 port map(XO0 => XO1, A0 => v114, OE => OE);
    vv113: XTRI1 port map(XO0 => XO2, A0 => v124, OE => OE);
    vv114: XTRI1 port map(XO0 => XO3, A0 => v134, OE => OE);
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT24E is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT24E;

architecture LATTICE_ARCH of ODT24E is
    signal v108, v118, v128, v138: std_logic;

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
      
    component XDFF2E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF2E use entity LAT_VHD.XDFF2E(LATTICE_ARCH);

begin
    v100: XTRI1 port map(XO0 => XO0, A0 => v108, OE => OE);
    v101: XTRI1 port map(XO0 => XO1, A0 => v118, OE => OE);
    v102: XTRI1 port map(XO0 => XO2, A0 => v128, OE => OE);
    v103: XTRI1 port map(XO0 => XO3, A0 => v138, OE => OE);

    v110: XDFF2E port map(Q0 => v108, D0 => D0, CLK => CLK, CD => CD, EN => EN);
    v111: XDFF2E port map(Q0 => v118, D0 => D1, CLK => CLK, CD => CD, EN => EN);
    v112: XDFF2E port map(Q0 => v128, D0 => D2, CLK => CLK, CD => CD, EN => EN);
    v113: XDFF2E port map(Q0 => v138, D0 => D3, CLK => CLK, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT31 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         OE: IN std_logic);
end ODT31;

architecture LATTICE_ARCH of ODT31 is
    signal v104: std_logic;
    
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v107: XDFF3
        port map(Q0 => v104,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD);
    
    v108: XTRI1
        port map(XO0 => XO0,
                 A0 => v104,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT31E is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic;
         OE: IN std_logic);
end ODT31E;

architecture LATTICE_ARCH of ODT31E is
    signal v108: std_logic;
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);
    
begin
    v111: XTRI1
        port map(XO0 => XO0,
                 A0 => v108,
                 OE => OE);
    
    v112: XDFF3E
        port map(Q0 => v108,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT34 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         OE: IN std_logic);
end ODT34;

architecture LATTICE_ARCH of ODT34 is
    signal v104, v114, v124, v134: std_logic;
    
    component XDFF3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDFF3 use entity LAT_VHD.XDFF3(LATTICE_ARCH);

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin
    v100: XDFF3 port map(Q0 => v104, D0 => D0, CLK => CLK, SD => SD);
    v101: XDFF3 port map(Q0 => v114, D0 => D1, CLK => CLK, SD => SD);
    v102: XDFF3 port map(Q0 => v124, D0 => D2, CLK => CLK, SD => SD);
    v103: XDFF3 port map(Q0 => v134, D0 => D3, CLK => CLK, SD => SD);

    v110: XTRI1 port map(XO0 => XO0, A0 => v104, OE => OE);
    v111: XTRI1 port map(XO0 => XO1, A0 => v114, OE => OE);
    v112: XTRI1 port map(XO0 => XO2, A0 => v124, OE => OE);
    v113: XTRI1 port map(XO0 => XO3, A0 => v134, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT34E is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end ODT34E;

architecture LATTICE_ARCH of ODT34E is
    signal v108, v118, v128, v138 : std_logic;

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
       
    component XDFF3E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF3E use entity LAT_VHD.XDFF3E(LATTICE_ARCH);

begin

    v100: XTRI1 port map(XO0 => XO0, A0 => v108, OE => OE);
    v101: XTRI1 port map(XO0 => XO1, A0 => v118, OE => OE);
    v102: XTRI1 port map(XO0 => XO2, A0 => v128, OE => OE);
    v103: XTRI1 port map(XO0 => XO3, A0 => v138, OE => OE);

    v110: XDFF3E port map(Q0 => v108, D0 => D0, CLK => CLK, SD => SD, EN => EN);
    v111: XDFF3E port map(Q0 => v118, D0 => D1, CLK => CLK, SD => SD, EN => EN);
    v112: XDFF3E port map(Q0 => v128, D0 => D2, CLK => CLK, SD => SD, EN => EN);
    v113: XDFF3E port map(Q0 => v138, D0 => D3, CLK => CLK, SD => SD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT41 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT41;

architecture LATTICE_ARCH of ODT41 is
    signal v101: std_logic;
    
    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v104: XDFF4
        port map(Q0 => v101,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v105: XTRI1
        port map(XO0 => XO0,
                 A0 => v101,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT41E is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         CLK: IN std_logic;
         EN: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT41E;

architecture LATTICE_ARCH of ODT41E is
    signal v105: std_logic;
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);
    
begin
    v108: XTRI1
        port map(XO0 => XO0,
                 A0 => v105,
                 OE => OE);
    
    v109: XDFF4E
        port map(Q0 => v105,
                 D0 => D0,
                 CLK => CLK,
                 SD => SD,
                 CD => CD,
                 EN => EN);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT44 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end ODT44;

architecture LATTICE_ARCH of ODT44 is
    signal v101, v111, v121, v131: std_logic;

    component XDFF4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDFF4 use entity LAT_VHD.XDFF4(LATTICE_ARCH);

    component XTRI1
    port(XO0: OUT std_logic;
         A0: IN std_logic;
         OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    vv100: XDFF4 port map(Q0 => v101, D0 => D0, CLK => CLK, SD => SD, CD => CD);
    vv101: XDFF4 port map(Q0 => v111, D0 => D1, CLK => CLK, SD => SD, CD => CD);
    vv102: XDFF4 port map(Q0 => v121, D0 => D2, CLK => CLK, SD => SD, CD => CD);
    vv103: XDFF4 port map(Q0 => v131, D0 => D3, CLK => CLK, SD => SD, CD => CD);

    vv110: XTRI1 port map(XO0 => XO0, A0 => v101, OE => OE);
    vv111: XTRI1 port map(XO0 => XO1, A0 => v111, OE => OE);
    vv112: XTRI1 port map(XO0 => XO2, A0 => v121, OE => OE);
    vv113: XTRI1 port map(XO0 => XO3, A0 => v131, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity ODT44E is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         EN: IN std_logic;
         OE: IN std_logic);
end ODT44E;

architecture LATTICE_ARCH of ODT44E is
    signal v105, v115, v125, v135: std_logic;

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
     
    component XDFF4E
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic;
             EN: IN std_logic);
    end component;
    for all : XDFF4E use entity LAT_VHD.XDFF4E(LATTICE_ARCH);

begin

    v100: XTRI1 port map(XO0 => XO0, A0 => v105, OE => OE);
    v101: XTRI1 port map(XO0 => XO1, A0 => v115, OE => OE);
    v102: XTRI1 port map(XO0 => XO2, A0 => v125, OE => OE);
    v103: XTRI1 port map(XO0 => XO3, A0 => v135, OE => OE);

    v110: XDFF4E port map(Q0 => v105, D0 => D0, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v111: XDFF4E port map(Q0 => v115, D0 => D1, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v112: XDFF4E port map(Q0 => v125, D0 => D2, CLK => CLK, SD => SD, CD => CD, EN => EN);
    v113: XDFF4E port map(Q0 => v135, D0 => D3, CLK => CLK, SD => SD, CD => CD, EN => EN);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL11 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic);
end OL11;

architecture LATTICE_ARCH of OL11 is
    
    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);
    
begin
    v101: XDL1
        port map(Q0 => XQ0,
                 D0 => D0,
                 G => G);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL14 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic);
end OL14;

architecture LATTICE_ARCH of OL14 is

    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);

begin
    v100: XDL1 port map(Q0 => XQ0, D0 => D0, G => G);
    v101: XDL1 port map(Q0 => XQ1, D0 => D1, G => G);
    v102: XDL1 port map(Q0 => XQ2, D0 => D2, G => G);
    v103: XDL1 port map(Q0 => XQ3, D0 => D3, G => G);
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL21 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic);
end OL21;

architecture LATTICE_ARCH of OL21 is
    signal v100: std_logic;
    
    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
begin
    v103: XDL1
        port map(Q0 => XQ0,
                 D0 => D0,
                 G => v100);
    
    v104: INV
        port map(ZN0 => v100,
                 A0 => G);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL24 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic);
end OL24;

architecture LATTICE_ARCH of OL24 is
    signal v100: std_logic;

    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all: XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);

begin

    vv100: XDL1 port map(Q0 => XQ0, D0 => D0, G => v100);
    vv101: XDL1 port map(Q0 => XQ1, D0 => D1, G => v100);
    vv102: XDL1 port map(Q0 => XQ2, D0 => D2, G => v100);
    vv103: XDL1 port map(Q0 => XQ3, D0 => D3, G => v100);

    vv110: INV port map(ZN0 => v100, A0 => G);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL31 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic);
end OL31;

architecture LATTICE_ARCH of OL31 is
    
    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);
    
begin
    v104: XDL2
        port map(Q0 => XQ0,
                 D0 => D0,
                 G => G,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL34 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic);
end OL34;

architecture LATTICE_ARCH of OL34 is

    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);

begin

    v100: XDL2 port map(Q0 => XQ0, D0 => D0, G => G, CD => CD);
    v101: XDL2 port map(Q0 => XQ1, D0 => D1, G => G, CD => CD);
    v102: XDL2 port map(Q0 => XQ2, D0 => D2, G => G, CD => CD);
    v103: XDL2 port map(Q0 => XQ3, D0 => D3, G => G, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL41 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic);
end OL41;

architecture LATTICE_ARCH of OL41 is
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);
    
begin
    v104: XDL3
        port map(Q0 => XQ0,
                 D0 => D0,
                 G => G,
                 SD => SD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL44 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic);
end OL44;

architecture LATTICE_ARCH of OL44 is
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all: XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);

begin

    v100: XDL3 port map(Q0 => XQ0, D0 => D0, G => G, SD => SD);
    v101: XDL3 port map(Q0 => XQ1, D0 => D1, G => G, SD => SD);
    v102: XDL3 port map(Q0 => XQ2, D0 => D2, G => G, SD => SD);
    v103: XDL3 port map(Q0 => XQ3, D0 => D3, G => G, SD => SD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL51 is
    port(XQ0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic);
end OL51;

architecture LATTICE_ARCH of OL51 is
    
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
    
begin
    v102: XDL4
        port map(Q0 => XQ0,
                 D0 => D0,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OL54 is
    port(XQ0: OUT std_logic;
         XQ1: OUT std_logic;
         XQ2: OUT std_logic;
         XQ3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic);
end OL54;

architecture LATTICE_ARCH of OL54 is

    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
							   
begin

    v100: XDL4 port map(Q0 => XQ0, D0 => D0, G => G, SD => SD, CD => CD);
    v101: XDL4 port map(Q0 => XQ1, D0 => D1, G => G, SD => SD, CD => CD);
    v102: XDL4 port map(Q0 => XQ2, D0 => D2, G => G, SD => SD, CD => CD);
    v103: XDL4 port map(Q0 => XQ3, D0 => D3, G => G, SD => SD, CD => CD);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT11 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end OLT11;

architecture LATTICE_ARCH of OLT11 is
    signal v101: std_logic;
    
    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all : XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v104: XDL1
        port map(Q0 => v101,
                 D0 => D0,
                 G => G);
    
    v105: XTRI1
        port map(XO0 => XO0,
                 A0 => v101,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT14 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         OE: IN std_logic);
end OLT14;

architecture LATTICE_ARCH of OLT14 is
    signal v101, v111, v121, v131: std_logic;
    
    component XDL1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic);
    end component;
    for all : XDL1 use entity LAT_VHD.XDL1(LATTICE_ARCH);
 
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    vv100: XDL1 port map(Q0 => v101, D0 => D0, G => G);
    vv101: XDL1 port map(Q0 => v111, D0 => D1, G => G);
    vv102: XDL1 port map(Q0 => v121, D0 => D2, G => G);
    vv103: XDL1 port map(Q0 => v131, D0 => D3, G => G);

    vv110: XTRI1 port map(XO0 => XO0, A0 => v101, OE => OE);
    vv111: XTRI1 port map(XO0 => XO1, A0 => v111, OE => OE);
    vv112: XTRI1 port map(XO0 => XO2, A0 => v121, OE => OE);
    vv113: XTRI1 port map(XO0 => XO3, A0 => v131, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT21 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end OLT21;

architecture LATTICE_ARCH of OLT21 is
    signal v104: std_logic;
    
    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v107: XDL2
        port map(Q0 => v104,
                 D0 => D0,
                 G => G,
                 CD => CD);
    
    v108: XTRI1
        port map(XO0 => XO0,
                 A0 => v104,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT24 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end OLT24;

architecture LATTICE_ARCH of OLT24 is
    signal v104, v114, v124, v134: std_logic;

    component XDL2
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL2 use entity LAT_VHD.XDL2(LATTICE_ARCH);
     
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    v100: XDL2 port map(Q0 => v104, D0 => D0, G => G, CD => CD);
    v101: XDL2 port map(Q0 => v114, D0 => D1, G => G, CD => CD);
    v102: XDL2 port map(Q0 => v124, D0 => D2, G => G, CD => CD);
    v103: XDL2 port map(Q0 => v134, D0 => D3, G => G, CD => CD);

    v110: XTRI1 port map(XO0 => XO0, A0 => v104, OE => OE);
    v111: XTRI1 port map(XO0 => XO1, A0 => v114, OE => OE);
    v112: XTRI1 port map(XO0 => XO2, A0 => v124, OE => OE);
    v113: XTRI1 port map(XO0 => XO3, A0 => v134, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT31 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic;
         OE: IN std_logic);
end OLT31;

architecture LATTICE_ARCH of OLT31 is
    signal v104: std_logic;
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v107: XDL3
        port map(Q0 => v104,
                 D0 => D0,
                 G => G,
                 SD => SD);
    
    v108: XTRI1
        port map(XO0 => XO0,
                 A0 => v104,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT34 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic;
         OE: IN std_logic);
end OLT34;

architecture LATTICE_ARCH of OLT34 is
    signal v104, v114, v124, v134: std_logic;
    
    component XDL3
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic);
    end component;
    for all : XDL3 use entity LAT_VHD.XDL3(LATTICE_ARCH);

    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    v100: XDL3 port map(Q0 => v104, D0 => D0, G => G, SD => SD);
    v101: XDL3 port map(Q0 => v114, D0 => D1, G => G, SD => SD);
    v102: XDL3 port map(Q0 => v124, D0 => D2, G => G, SD => SD);
    v103: XDL3 port map(Q0 => v134, D0 => D3, G => G, SD => SD);

    v110: XTRI1 port map(XO0 => XO0, A0 => v104, OE => OE);
    v111: XTRI1 port map(XO0 => XO1, A0 => v114, OE => OE);
    v112: XTRI1 port map(XO0 => XO2, A0 => v124, OE => OE);
    v113: XTRI1 port map(XO0 => XO3, A0 => v134, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT41 is
    port(XO0: OUT std_logic;
         D0: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end OLT41;

architecture LATTICE_ARCH of OLT41 is
    signal v102: std_logic;
    
    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
    
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);
    
begin
    v105: XDL4
        port map(Q0 => v102,
                 D0 => D0,
                 G => G,
                 SD => SD,
                 CD => CD);
    
    v106: XTRI1
        port map(XO0 => XO0,
                 A0 => v102,
                 OE => OE);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity OLT44 is
    port(XO0: OUT std_logic;
         XO1: OUT std_logic;
         XO2: OUT std_logic;
         XO3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         G: IN std_logic;
         SD: IN std_logic;
         CD: IN std_logic;
         OE: IN std_logic);
end OLT44;

architecture LATTICE_ARCH of OLT44 is
    signal v102, v112, v122, v132: std_logic;

    component XDL4
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             G: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all : XDL4 use entity LAT_VHD.XDL4(LATTICE_ARCH);
  
    component XTRI1
        port(XO0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all : XTRI1 use entity LAT_VHD.XTRI1(LATTICE_ARCH);

begin

    vv100: XDL4 port map(Q0 => v102, D0 => D0, G => G, SD => SD, CD => CD);
    vv101: XDL4 port map(Q0 => v112, D0 => D1, G => G, SD => SD, CD => CD);
    vv102: XDL4 port map(Q0 => v122, D0 => D2, G => G, SD => SD, CD => CD);
    vv103: XDL4 port map(Q0 => v132, D0 => D3, G => G, SD => SD, CD => CD);

    vv110: XTRI1 port map(XO0 => XO0, A0 => v102, OE => OE);
    vv111: XTRI1 port map(XO0 => XO1, A0 => v112, OE => OE);
    vv112: XTRI1 port map(XO0 => XO2, A0 => v122, OE => OE);
    vv113: XTRI1 port map(XO0 => XO3, A0 => v132, OE => OE);

end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity SRR51 is
    port(Q0: OUT std_logic;
         D0: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic);
end SRR51;

architecture LATTICE_ARCH of SRR51 is
    signal v101: std_logic;
    signal v102: std_logic;
    signal v106: std_logic;
    signal v100: std_logic;
    signal v103: std_logic;
    signal v104: std_logic;
    signal v105: std_logic;
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all: AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component OR3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: OR3 use entity LAT_VHD.OR3(LATTICE_ARCH);
    
begin
    v115: INV
        port map(ZN0 => v105,
                 A0 => EN);
    
    v116: INV
        port map(ZN0 => v100,
                 A0 => LD);
    
    v117: AND2
        port map(Z0 => v101,
                 A0 => LD,
                 A1 => D0);
    
    v118: AND3
        port map(Z0 => v103,
                 A0 => EN,
                 A1 => v100,
                 A2 => CAI);
    
    v119: BUF
        port map(Z0 => Q0,
                 A0 => v106);
    
    v120: AND3
        port map(Z0 => v102,
                 A0 => v106,
                 A1 => v100,
                 A2 => v105);
    
    v121: FDE1
        port map(Q0 => v106,
                 D0 => v104,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v122: OR3
        port map(Z0 => v104,
                 A0 => v102,
                 A1 => v103,
                 A2 => v101);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity SRR54 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic);
end SRR54;

architecture LATTICE_ARCH of SRR54 is
    signal v107: std_logic;
    signal v109: std_logic;
    signal v108: std_logic;
    signal v101, v111, v121, v131: std_logic;
    signal v102, v112, v122, v132: std_logic;
    signal v106, v116, v126, v136: std_logic;
    signal v100: std_logic;
    signal v103, v113, v123, v133: std_logic;
    signal v104, v114, v124, v134: std_logic;
    signal v105: std_logic;
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
   
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all: AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);

    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);

    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
   
    component OR3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: OR3 use entity LAT_VHD.OR3(LATTICE_ARCH);

begin
    
    vv100: BUF port map(Z0 => Q0, A0 => v107);
    vv101: BUF port map(Z0 => Q1, A0 => v108);
    vv102: BUF port map(Z0 => Q2, A0 => v109);
    
    vv103: INV port map(ZN0 => v105, A0 => EN);
    vv104: INV port map(ZN0 => v100, A0 => LD);

    vv110: AND2 port map(Z0 => v101, A0 => LD, A1 => D0);
    vv111: AND2 port map(Z0 => v111, A0 => LD, A1 => D1);
    vv112: AND2 port map(Z0 => v121, A0 => LD, A1 => D2);
    vv113: AND2 port map(Z0 => v131, A0 => LD, A1 => D3);

    vv120: AND3 port map(Z0 => v103, A0 => EN, A1 => v100, A2 => CAI);
    vv121: AND3 port map(Z0 => v113, A0 => EN, A1 => v100, A2 => V107);
    vv122: AND3 port map(Z0 => v123, A0 => EN, A1 => v100, A2 => V108);
    vv123: AND3 port map(Z0 => v133, A0 => EN, A1 => v100, A2 => V109);

    vv130: BUF port map(Z0 => v107, A0 => v106);
    vv131: BUF port map(Z0 => v108, A0 => v116);
    vv132: BUF port map(Z0 => v109, A0 => v126);
    vv133: BUF port map(Z0 => Q3, A0 => v136);

    vv140: AND3 port map(Z0 => v102, A0 => v106, A1 => v100, A2 => v105);
    vv141: AND3 port map(Z0 => v112, A0 => v116, A1 => v100, A2 => v105);
    vv142: AND3 port map(Z0 => v122, A0 => v126, A1 => v100, A2 => v105);
    vv143: AND3 port map(Z0 => v132, A0 => v136, A1 => v100, A2 => v105);

    vv150: FDE1 port map(Q0 => v106, D0 => v104, CLK => CLK, SD => SD, CD => CD);
    vv151: FDE1 port map(Q0 => v116, D0 => v114, CLK => CLK, SD => SD, CD => CD);
    vv152: FDE1 port map(Q0 => v126, D0 => v124, CLK => CLK, SD => SD, CD => CD);
    vv153: FDE1 port map(Q0 => v136, D0 => v134, CLK => CLK, SD => SD, CD => CD);

    vv160: OR3 port map(Z0 => v104, A0 => v102, A1 => v103, A2 => v101);
    vv161: OR3 port map(Z0 => v114, A0 => v112, A1 => v113, A2 => v111);
    vv162: OR3 port map(Z0 => v124, A0 => v122, A1 => v123, A2 => v121);
    vv163: OR3 port map(Z0 => v134, A0 => v132, A1 => v133, A2 => v131);
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity SRR58 is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAI: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         CD: IN std_logic);
end SRR58;

architecture LATTICE_ARCH of SRR58 is
    signal v107, v117, v127, v137, v147, v157, v167: std_logic;
    signal v101, v111, v121, v131, v141, v151, v161, v171: std_logic;
    signal v102, v112, v122, v132, v142, v152, v162, v172: std_logic;
    signal v106, v116, v126, v136, v146, v156, v166, v176: std_logic;
    signal v100: std_logic;
    signal v103, v113, v123, v133, v143, v153, v163, v173: std_logic;
    signal v104, v114, v124, v134, v144, v154, v164, v174: std_logic;
    signal v105: std_logic;
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: BUF use entity LAT_VHD.BUF(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
   
    component AND2
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic);
    end component;
    for all: AND2 use entity LAT_VHD.AND2(LATTICE_ARCH);

    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);

    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
   
    component OR3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: OR3 use entity LAT_VHD.OR3(LATTICE_ARCH);

begin

    vv100: BUF port map(Z0 => Q0, A0 => v107);
    vv101: BUF port map(Z0 => Q1, A0 => v117);
    vv102: BUF port map(Z0 => Q2, A0 => v127);
    vv103: BUF port map(Z0 => Q3, A0 => v137);
    vv104: BUF port map(Z0 => Q4, A0 => v147);
    vv105: BUF port map(Z0 => Q5, A0 => v157);
    vv106: BUF port map(Z0 => Q6, A0 => v167);
    
    vv107: INV port map(ZN0 => v105, A0 => EN);
    vv108: INV port map(ZN0 => v100, A0 => LD);

    vv110: AND2 port map(Z0 => v101, A0 => LD, A1 => D0);
    vv111: AND2 port map(Z0 => v111, A0 => LD, A1 => D1);
    vv112: AND2 port map(Z0 => v121, A0 => LD, A1 => D2);
    vv113: AND2 port map(Z0 => v131, A0 => LD, A1 => D3);
    vv114: AND2 port map(Z0 => v141, A0 => LD, A1 => D4);
    vv115: AND2 port map(Z0 => v151, A0 => LD, A1 => D5);
    vv116: AND2 port map(Z0 => v161, A0 => LD, A1 => D6);
    vv117: AND2 port map(Z0 => v171, A0 => LD, A1 => D7);

    vv120: AND3 port map(Z0 => v103, A0 => EN, A1 => v100, A2 => CAI);
    vv121: AND3 port map(Z0 => v113, A0 => EN, A1 => v100, A2 => V107);
    vv122: AND3 port map(Z0 => v123, A0 => EN, A1 => v100, A2 => V117);
    vv123: AND3 port map(Z0 => v133, A0 => EN, A1 => v100, A2 => V127);
    vv124: AND3 port map(Z0 => v143, A0 => EN, A1 => v100, A2 => V137);
    vv125: AND3 port map(Z0 => v153, A0 => EN, A1 => v100, A2 => V147);
    vv126: AND3 port map(Z0 => v163, A0 => EN, A1 => v100, A2 => V157);
    vv127: AND3 port map(Z0 => v173, A0 => EN, A1 => v100, A2 => V167);

    vv130: BUF port map(Z0 => v107, A0 => v106);
    vv131: BUF port map(Z0 => v117, A0 => v116);
    vv132: BUF port map(Z0 => v127, A0 => v126);
    vv133: BUF port map(Z0 => v137, A0 => v136);
    vv134: BUF port map(Z0 => v147, A0 => v146);
    vv135: BUF port map(Z0 => v157, A0 => v156);
    vv136: BUF port map(Z0 => v167, A0 => v166);
    vv137: BUF port map(Z0 => Q7, A0 => v176);

    vv140: AND3 port map(Z0 => v102, A0 => v106, A1 => v100, A2 => v105);
    vv141: AND3 port map(Z0 => v112, A0 => v116, A1 => v100, A2 => v105);
    vv142: AND3 port map(Z0 => v122, A0 => v126, A1 => v100, A2 => v105);
    vv143: AND3 port map(Z0 => v132, A0 => v136, A1 => v100, A2 => v105);
    vv144: AND3 port map(Z0 => v142, A0 => v146, A1 => v100, A2 => v105);
    vv145: AND3 port map(Z0 => v152, A0 => v156, A1 => v100, A2 => v105);
    vv146: AND3 port map(Z0 => v162, A0 => v166, A1 => v100, A2 => v105);
    vv147: AND3 port map(Z0 => v172, A0 => v176, A1 => v100, A2 => v105);

    vv150: FDE1 port map(Q0 => v106, D0 => v104, CLK => CLK, SD => SD, CD => CD);
    vv151: FDE1 port map(Q0 => v116, D0 => v114, CLK => CLK, SD => SD, CD => CD);
    vv152: FDE1 port map(Q0 => v126, D0 => v124, CLK => CLK, SD => SD, CD => CD);
    vv153: FDE1 port map(Q0 => v136, D0 => v134, CLK => CLK, SD => SD, CD => CD);
    vv154: FDE1 port map(Q0 => v146, D0 => v144, CLK => CLK, SD => SD, CD => CD);
    vv155: FDE1 port map(Q0 => v156, D0 => v154, CLK => CLK, SD => SD, CD => CD);
    vv156: FDE1 port map(Q0 => v166, D0 => v164, CLK => CLK, SD => SD, CD => CD);
    vv157: FDE1 port map(Q0 => v176, D0 => v174, CLK => CLK, SD => SD, CD => CD);

    vv160: OR3 port map(Z0 => v104, A0 => v102, A1 => v103, A2 => v101);
    vv161: OR3 port map(Z0 => v114, A0 => v112, A1 => v113, A2 => v111);
    vv162: OR3 port map(Z0 => v124, A0 => v122, A1 => v123, A2 => v121);
    vv163: OR3 port map(Z0 => v134, A0 => v132, A1 => v133, A2 => v131);
    vv164: OR3 port map(Z0 => v144, A0 => v142, A1 => v143, A2 => v141);
    vv165: OR3 port map(Z0 => v154, A0 => v152, A1 => v153, A2 => v151);
    vv166: OR3 port map(Z0 => v164, A0 => v162, A1 => v163, A2 => v161);
    vv167: OR3 port map(Z0 => v174, A0 => v172, A1 => v173, A2 => v171);
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity SRRL1S is
    port(Q0: OUT std_logic;
         D0: IN std_logic;
         CAIR: IN std_logic;
         CAIL: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         PS: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         RL: IN std_logic;
         CD: IN std_logic;
         CS: IN std_logic);
end SRRL1S;

architecture LATTICE_ARCH of SRRL1S is
    signal v100: std_logic;
    signal v103: std_logic;
    signal v104: std_logic;
    signal v101: std_logic;
    signal v107: std_logic;
    signal v105: std_logic;
    signal v102: std_logic;
    signal v106: std_logic;
    signal v109: std_logic;
    signal v108: std_logic;
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all: AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
    
    component OR5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all: OR5 use entity LAT_VHD.OR5(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
    
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);
    
    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
    
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all: AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);
    
begin
    v121: AND4
        port map(Z0 => v101,
                 A0 => v107,
                 A1 => v106,
                 A2 => v108,
                 A3 => v109);
    
    v122: OR5
        port map(Z0 => v105,
                 A0 => v101,
                 A1 => v102,
                 A2 => v103,
                 A3 => v104,
                 A4 => PS);
    
    v123: INV
        port map(ZN0 => v100,
                 A0 => RL);
    
    v124: INV
        port map(ZN0 => v109,
                 A0 => CS);
    
    v125: INV
        port map(ZN0 => v106,
                 A0 => LD);
    
    v126: INV
        port map(ZN0 => v108,
                 A0 => EN);
    
    v127: BUF
        port map(Z0 => Q0,
                 A0 => v107);
    
    v128: AND3
        port map(Z0 => v104,
                 A0 => LD,
                 A1 => v109,
                 A2 => D0);
    
    v129: FDE1
        port map(Q0 => v107,
                 D0 => v105,
                 CLK => CLK,
                 SD => SD,
                 CD => CD);
    
    v130: AND5
        port map(Z0 => v102,
                 A0 => EN,
                 A1 => v106,
                 A2 => v109,
                 A3 => RL,
                 A4 => CAIR);
    
    v131: AND5
        port map(Z0 => v103,
                 A0 => EN,
                 A1 => v106,
                 A2 => v109,
                 A3 => v100,
                 A4 => CAIL);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity SRRL4S is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         CAIR: IN std_logic;
         CAIL: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         PS: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         RL: IN std_logic;
         CD: IN std_logic;
         CS: IN std_logic);
end SRRL4S;

architecture LATTICE_ARCH of SRRL4S is
    signal v100: std_logic;
    signal v106: std_logic;
    signal v108: std_logic;
    signal v109: std_logic;
    signal v101, v111, v121, v131: std_logic;
    signal v102, v112, v122, v132: std_logic;
    signal v103, v113, v123, v133: std_logic;
    signal v104, v114, v124, v134: std_logic;
    signal v105, v115, v125, v135: std_logic;
    signal v107, v117, v127, v137: std_logic;
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all: AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
   
    component OR5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all: OR5 use entity LAT_VHD.OR5(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
   
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
        
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);

    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
   
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all: AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);

begin
    
    vv100: INV port map(ZN0 => v100, A0 => RL);
    vv101: INV port map(ZN0 => v109, A0 => CS);
    vv102: INV port map(ZN0 => v106, A0 => LD);
    vv103: INV port map(ZN0 => v108, A0 => EN);

    vv110: AND4 port map(Z0 => v101, A0 => v107, A1 => v106, A2 => v108, A3 => v109);
    vv111: AND4 port map(Z0 => v111, A0 => v117, A1 => v106, A2 => v108, A3 => v109);
    vv112: AND4 port map(Z0 => v121, A0 => v127, A1 => v106, A2 => v108, A3 => v109);
    vv113: AND4 port map(Z0 => v131, A0 => v137, A1 => v106, A2 => v108, A3 => v109);

    vv120: OR5 port map(Z0 => v105, A0 => v101, A1 => v102, A2 => v103, A3 => v104, A4 => PS);
    vv121: OR5 port map(Z0 => v115, A0 => v111, A1 => v112, A2 => v113, A3 => v114, A4 => PS);
    vv122: OR5 port map(Z0 => v125, A0 => v121, A1 => v122, A2 => v123, A3 => v124, A4 => PS);
    vv123: OR5 port map(Z0 => v135, A0 => v131, A1 => v132, A2 => v133, A3 => v134, A4 => PS);

    vv130: BUF port map(Z0 => Q0, A0 => v107);
    vv131: BUF port map(Z0 => Q1, A0 => v117);
    vv132: BUF port map(Z0 => Q2, A0 => v127);
    vv133: BUF port map(Z0 => Q3, A0 => v137);

    vv140: AND3 port map(Z0 => v104, A0 => LD, A1 => v109, A2 => D0);
    vv141: AND3 port map(Z0 => v114, A0 => LD, A1 => v109, A2 => D1);
    vv142: AND3 port map(Z0 => v124, A0 => LD, A1 => v109, A2 => D2);
    vv143: AND3 port map(Z0 => v134, A0 => LD, A1 => v109, A2 => D3);

    vv150: FDE1 port map(Q0 => v107, D0 => v105, CLK => CLK, SD => SD, CD => CD);
    vv151: FDE1 port map(Q0 => v117, D0 => v115, CLK => CLK, SD => SD, CD => CD);
    vv152: FDE1 port map(Q0 => v127, D0 => v125, CLK => CLK, SD => SD, CD => CD);
    vv153: FDE1 port map(Q0 => v137, D0 => v135, CLK => CLK, SD => SD, CD => CD);

    vv160: AND5 port map(Z0 => v102, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => CAIR);
    vv161: AND5 port map(Z0 => v112, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V107);
    vv162: AND5 port map(Z0 => v122, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V117);
    vv163: AND5 port map(Z0 => v132, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V127);

    vv170: AND5 port map(Z0 => v103, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V117);
    vv171: AND5 port map(Z0 => v113, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V127);
    vv172: AND5 port map(Z0 => v123, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V137);
    vv173: AND5 port map(Z0 => v133, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => CAIL);
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity SRRL8S is
    port(Q0: OUT std_logic;
         Q1: OUT std_logic;
         Q2: OUT std_logic;
         Q3: OUT std_logic;
         Q4: OUT std_logic;
         Q5: OUT std_logic;
         Q6: OUT std_logic;
         Q7: OUT std_logic;
         D0: IN std_logic;
         D1: IN std_logic;
         D2: IN std_logic;
         D3: IN std_logic;
         D4: IN std_logic;
         D5: IN std_logic;
         D6: IN std_logic;
         D7: IN std_logic;
         CAIR: IN std_logic;
         CAIL: IN std_logic;
         CLK: IN std_logic;
         SD: IN std_logic;
         PS: IN std_logic;
         LD: IN std_logic;
         EN: IN std_logic;
         RL: IN std_logic;
         CD: IN std_logic;
         CS: IN std_logic);
end SRRL8S;

architecture LATTICE_ARCH of SRRL8S is
    signal v100: std_logic;
    signal v106: std_logic;
    signal v108: std_logic;
    signal v109: std_logic;
    signal v101, v111, v121, v131, v141, v151, v161, v171: std_logic;
    signal v102, v112, v122, v132, v142, v152, v162, v172: std_logic;
    signal v103, v113, v123, v133, v143, v153, v163, v173: std_logic;
    signal v104, v114, v124, v134, v144, v154, v164, v174: std_logic;
    signal v105, v115, v125, v135, v145, v155, v165, v175: std_logic;
    signal v107, v117, v127, v137, v147, v157, v167, v177: std_logic;
    
    component AND4
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic);
    end component;
    for all: AND4 use entity LAT_VHD.AND4(LATTICE_ARCH);
   
    component OR5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all: OR5 use entity LAT_VHD.OR5(LATTICE_ARCH);

    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
   
    component BUF
        port(Z0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: BUF use entity LAT_VHD.BUF(LATTICE_ARCH);
        
    component AND3
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic);
    end component;
    for all: AND3 use entity LAT_VHD.AND3(LATTICE_ARCH);

    component FDE1
        port(Q0: OUT std_logic;
             D0: IN std_logic;
             CLK: IN std_logic;
             SD: IN std_logic;
             CD: IN std_logic);
    end component;
    for all: FDE1 use entity LAT_VHD.FDE1(LATTICE_ARCH);
   
    component AND5
        port(Z0: OUT std_logic;
             A0: IN std_logic;
             A1: IN std_logic;
             A2: IN std_logic;
             A3: IN std_logic;
             A4: IN std_logic);
    end component;
    for all: AND5 use entity LAT_VHD.AND5(LATTICE_ARCH);

begin
    
    vv100: INV port map(ZN0 => v100, A0 => RL);
    vv101: INV port map(ZN0 => v109, A0 => CS);
    vv102: INV port map(ZN0 => v106, A0 => LD);
    vv103: INV port map(ZN0 => v108, A0 => EN);

    vv110: AND4 port map(Z0 => v101, A0 => v107, A1 => v106, A2 => v108, A3 => v109);
    vv111: AND4 port map(Z0 => v111, A0 => v117, A1 => v106, A2 => v108, A3 => v109);
    vv112: AND4 port map(Z0 => v121, A0 => v127, A1 => v106, A2 => v108, A3 => v109);
    vv113: AND4 port map(Z0 => v131, A0 => v137, A1 => v106, A2 => v108, A3 => v109);
    vv114: AND4 port map(Z0 => v141, A0 => v147, A1 => v106, A2 => v108, A3 => v109);
    vv115: AND4 port map(Z0 => v151, A0 => v157, A1 => v106, A2 => v108, A3 => v109);
    vv116: AND4 port map(Z0 => v161, A0 => v167, A1 => v106, A2 => v108, A3 => v109);
    vv117: AND4 port map(Z0 => v171, A0 => v177, A1 => v106, A2 => v108, A3 => v109);

    vv120: OR5 port map(Z0 => v105, A0 => v101, A1 => v102, A2 => v103, A3 => v104, A4 => PS);
    vv121: OR5 port map(Z0 => v115, A0 => v111, A1 => v112, A2 => v113, A3 => v114, A4 => PS);
    vv122: OR5 port map(Z0 => v125, A0 => v121, A1 => v122, A2 => v123, A3 => v124, A4 => PS);
    vv123: OR5 port map(Z0 => v135, A0 => v131, A1 => v132, A2 => v133, A3 => v134, A4 => PS);
    vv124: OR5 port map(Z0 => v145, A0 => v141, A1 => v142, A2 => v143, A3 => v144, A4 => PS);
    vv125: OR5 port map(Z0 => v155, A0 => v151, A1 => v152, A2 => v153, A3 => v154, A4 => PS);
    vv126: OR5 port map(Z0 => v165, A0 => v161, A1 => v162, A2 => v163, A3 => v164, A4 => PS);
    vv127: OR5 port map(Z0 => v175, A0 => v171, A1 => v172, A2 => v173, A3 => v174, A4 => PS);

    vv130: BUF port map(Z0 => Q0, A0 => v107);
    vv131: BUF port map(Z0 => Q1, A0 => v117);
    vv132: BUF port map(Z0 => Q2, A0 => v127);
    vv133: BUF port map(Z0 => Q3, A0 => v137);
    vv134: BUF port map(Z0 => Q4, A0 => v147);
    vv135: BUF port map(Z0 => Q5, A0 => v157);
    vv136: BUF port map(Z0 => Q6, A0 => v167);
    vv137: BUF port map(Z0 => Q7, A0 => v177);

    vv140: AND3 port map(Z0 => v104, A0 => LD, A1 => v109, A2 => D0);
    vv141: AND3 port map(Z0 => v114, A0 => LD, A1 => v109, A2 => D1);
    vv142: AND3 port map(Z0 => v124, A0 => LD, A1 => v109, A2 => D2);
    vv143: AND3 port map(Z0 => v134, A0 => LD, A1 => v109, A2 => D3);
    vv144: AND3 port map(Z0 => v144, A0 => LD, A1 => v109, A2 => D4);
    vv145: AND3 port map(Z0 => v154, A0 => LD, A1 => v109, A2 => D5);
    vv146: AND3 port map(Z0 => v164, A0 => LD, A1 => v109, A2 => D6);
    vv147: AND3 port map(Z0 => v174, A0 => LD, A1 => v109, A2 => D7);

    vv150: FDE1 port map(Q0 => v107, D0 => v105, CLK => CLK, SD => SD, CD => CD);
    vv151: FDE1 port map(Q0 => v117, D0 => v115, CLK => CLK, SD => SD, CD => CD);
    vv152: FDE1 port map(Q0 => v127, D0 => v125, CLK => CLK, SD => SD, CD => CD);
    vv153: FDE1 port map(Q0 => v137, D0 => v135, CLK => CLK, SD => SD, CD => CD);
    vv154: FDE1 port map(Q0 => v147, D0 => v145, CLK => CLK, SD => SD, CD => CD);
    vv155: FDE1 port map(Q0 => v157, D0 => v155, CLK => CLK, SD => SD, CD => CD);
    vv156: FDE1 port map(Q0 => v167, D0 => v165, CLK => CLK, SD => SD, CD => CD);
    vv157: FDE1 port map(Q0 => v177, D0 => v175, CLK => CLK, SD => SD, CD => CD);

    vv160: AND5 port map(Z0 => v102, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => CAIR);
    vv161: AND5 port map(Z0 => v112, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V107);
    vv162: AND5 port map(Z0 => v122, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V117);
    vv163: AND5 port map(Z0 => v132, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V127);
    vv164: AND5 port map(Z0 => v142, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V137);
    vv165: AND5 port map(Z0 => v152, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V147);
    vv166: AND5 port map(Z0 => v162, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V157);
    vv167: AND5 port map(Z0 => v172, A0 => EN, A1 => v106, A2 => v109, A3 => RL, A4 => V167);

    vv170: AND5 port map(Z0 => v103, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V117);
    vv171: AND5 port map(Z0 => v113, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V127);
    vv172: AND5 port map(Z0 => v123, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V137);
    vv173: AND5 port map(Z0 => v133, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V147);
    vv174: AND5 port map(Z0 => v143, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V157);
    vv175: AND5 port map(Z0 => v153, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V167);
    vv176: AND5 port map(Z0 => v163, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => V177);
    vv177: AND5 port map(Z0 => v173, A0 => EN, A1 => v106, A2 => v109, A3 => v100, A4 => CAIL);
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity TCVRDC is
    port(A: INOUT std_logic;
         B: INOUT std_logic;
         ENA: IN std_logic;
         ENB: IN std_logic);
end TCVRDC;

architecture LATTICE_ARCH of TCVRDC is
    
    component IT11
        port(O0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);
    
begin
    v103: IT11
        port map(O0 => B,
                 A0 => A,
                 OE => ENA);
    
    v104: IT11
        port map(O0 => A,
                 A0 => B,
                 OE => ENB);
    
    
end LATTICE_ARCH;
Library IEEE; 
Library LAT_VHD;
Use IEEE.STD_LOGIC_1164.all;
Use LAT_VHD.VHD_PKG.all;

entity TCVRSC is
    port(A: INOUT std_logic;
         B: INOUT std_logic;
         EN: IN std_logic);
end TCVRSC;

architecture LATTICE_ARCH of TCVRSC is
    signal v101: std_logic;
    
    component IT11
        port(O0: OUT std_logic;
             A0: IN std_logic;
             OE: IN std_logic);
    end component;
    for all: IT11 use entity LAT_VHD.IT11(LATTICE_ARCH);
    
    component INV
        port(ZN0: OUT std_logic;
             A0: IN std_logic);
    end component;
    for all: INV use entity LAT_VHD.INV(LATTICE_ARCH);
    
begin
    v105: IT11
        port map(O0 => B,
                 A0 => A,
                 OE => EN);
    
    v106: INV
        port map(ZN0 => v101,
                 A0 => EN);
    
    v107: IT11
        port map(O0 => A,
                 A0 => B,
                 OE => v101);
    
    
end LATTICE_ARCH;
