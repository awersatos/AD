// --------------------------------------------------------------------
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// --------------------------------------------------------------------
// Copyright (c) 2005 by Lattice Semiconductor Corporation
// --------------------------------------------------------------------
//
//
//                     Lattice Semiconductor Corporation
//                     5555 NE Moore Court
//                     Hillsboro, OR 97214
//                     U.S.A.
//
//                     TEL: 1-800-Lattice  (USA and Canada)
//                          1-408-826-6000 (other locations)
//
//                     web: http://www.latticesemi.com/
//                     email: techsupport@latticesemi.com
//
// --------------------------------------------------------------------
//
// Simulation Library File for ORCA4
//
// $Header: /home/dmsys/pvcs/RCSMigTest/rcs/verilog/pkg/versclibs/data/orca4/RCS/ULIM.v,v 1.2 2005/05/19 19:02:19 pradeep Exp $ 
//
`timescale 1 ns / 1 ps

`celldefine

module ULIM (ADDR0, ADDR1, ADDR2, ADDR3, ADDR4, ADDR5, ADDR6, ADDR7, ADDR8, ADDR9, ADDR10,
             ADDR11, ADDR12, ADDR13, ADDR14, ADDR15, ADDR16, ADDR17, WDATA0, WDATA1, WDATA2,
             WDATA3, WDATA4, WDATA5, WDATA6, WDATA7, WDATA8, WDATA9, WDATA10, WDATA11,
             WDATA12, WDATA13, WDATA14, WDATA15, WDATA16, WDATA17, WDATA18, WDATA19, WDATA20,
             WDATA21, WDATA22, WDATA23, WDATA24, WDATA25, WDATA26, WDATA27, WDATA28, WDATA29,
             WDATA30, WDATA31, WDATA32, WDATA33, WDATA34, WDATA35, CLK, RESET, WRITE, READ,
             BURST, RDY, SIZE0, SIZE1, LOCK, IRQ, SRDATA0, SRDATA1, SRDATA2, SRDATA3,
             SRDATA4, SRDATA5, SRDATA6, SRDATA7, SRDATA8, SRDATA9, SRDATA10, SRDATA11, 
             SRDATA12, SRDATA13, SRDATA14, SRDATA15, SRDATA16, SRDATA17, SRDATA18,
             SRDATA19, SRDATA20, SRDATA21, SRDATA22, SRDATA23, SRDATA24, SRDATA25,
             SRDATA26, SRDATA27, SRDATA28, SRDATA29, SRDATA30, SRDATA31, SRDATA32,
             SRDATA33, SRDATA34, SRDATA35, SGRANTED, SACK, SRETRY, SERR,
             RDATA0, RDATA1, RDATA2, RDATA3, RDATA4, RDATA5, RDATA6, RDATA7, RDATA8,
             RDATA9, RDATA10, RDATA11, RDATA12, RDATA13, RDATA14, RDATA15, RDATA16, RDATA17,
             RDATA18, RDATA19, RDATA20, RDATA21, RDATA22, RDATA23, RDATA24, RDATA25, RDATA26,
             RDATA27, RDATA28, RDATA29, RDATA30, RDATA31, RDATA32, RDATA33, RDATA34, RDATA35,
             GRANTED, ACK, RETRY, ERR, SADDR0, SADDR1, SADDR2, SADDR3, SADDR4, SADDR5,
             SADDR6, SADDR7, SADDR8, SADDR9, SADDR10, SADDR11, SADDR12, SADDR13, SADDR14,
             SADDR15, SADDR16, SADDR17, SWDATA0, SWDATA1, SWDATA2, SWDATA3, SWDATA4, SWDATA5,
             SWDATA6, SWDATA7, SWDATA8, SWDATA9, SWDATA10, SWDATA11, SWDATA12, SWDATA13,
             SWDATA14, SWDATA15, SWDATA16, SWDATA17, SWDATA18, SWDATA19, SWDATA20,
             SWDATA21, SWDATA22, SWDATA23, SWDATA24, SWDATA25, SWDATA26, SWDATA27,
             SWDATA28, SWDATA29, SWDATA30, SWDATA31, SWDATA32, SWDATA33, SWDATA34, SWDATA35,
             SCLK, SRESET, SWRITE, SREAD, SBURST, SRDY, SSIZE0, SSIZE1, SLOCK, SIRQ);

input ADDR0, ADDR1, ADDR2, ADDR3, ADDR4, ADDR5, ADDR6, ADDR7, ADDR8, ADDR9, ADDR10;
input ADDR11, ADDR12, ADDR13, ADDR14, ADDR15, ADDR16, ADDR17, WDATA0, WDATA1, WDATA2;
input WDATA3, WDATA4, WDATA5, WDATA6, WDATA7, WDATA8, WDATA9, WDATA10, WDATA11;
input WDATA12, WDATA13, WDATA14, WDATA15, WDATA16, WDATA17, WDATA18, WDATA19, WDATA20;
input WDATA21, WDATA22, WDATA23, WDATA24, WDATA25, WDATA26, WDATA27, WDATA28, WDATA29;
input WDATA30, WDATA31, WDATA32, WDATA33, WDATA34, WDATA35, CLK, RESET, WRITE, READ;
input BURST, RDY, SIZE0, SIZE1, LOCK, IRQ, SRDATA0, SRDATA1, SRDATA2, SRDATA3;
input SRDATA4, SRDATA5, SRDATA6, SRDATA7, SRDATA8, SRDATA9, SRDATA10, SRDATA11;
input SRDATA12, SRDATA13, SRDATA14, SRDATA15, SRDATA16, SRDATA17, SRDATA18;
input SRDATA19, SRDATA20, SRDATA21, SRDATA22, SRDATA23, SRDATA24, SRDATA25;
input SRDATA26, SRDATA27, SRDATA28, SRDATA29, SRDATA30, SRDATA31, SRDATA32;
input SRDATA33, SRDATA34, SRDATA35, SGRANTED, SACK, SRETRY, SERR;

output RDATA0, RDATA1, RDATA2, RDATA3, RDATA4, RDATA5, RDATA6, RDATA7, RDATA8;
output RDATA9, RDATA10, RDATA11, RDATA12, RDATA13, RDATA14, RDATA15, RDATA16, RDATA17;
output RDATA18, RDATA19, RDATA20, RDATA21, RDATA22, RDATA23, RDATA24, RDATA25, RDATA26;
output RDATA27, RDATA28, RDATA29, RDATA30, RDATA31, RDATA32, RDATA33, RDATA34, RDATA35;
output GRANTED, ACK, RETRY, ERR, SADDR0, SADDR1, SADDR2, SADDR3, SADDR4, SADDR5;
output SADDR6, SADDR7, SADDR8, SADDR9, SADDR10, SADDR11, SADDR12, SADDR13, SADDR14;
output SADDR15, SADDR16, SADDR17, SWDATA0, SWDATA1, SWDATA2, SWDATA3, SWDATA4, SWDATA5;
output SWDATA6, SWDATA7, SWDATA8, SWDATA9, SWDATA10, SWDATA11, SWDATA12, SWDATA13;
output SWDATA14, SWDATA15, SWDATA16, SWDATA17, SWDATA18, SWDATA19, SWDATA20;
output SWDATA21, SWDATA22, SWDATA23, SWDATA24, SWDATA25, SWDATA26, SWDATA27;
output SWDATA28, SWDATA29, SWDATA30, SWDATA31, SWDATA32, SWDATA33, SWDATA34, SWDATA35;
output SCLK, SRESET, SWRITE, SREAD, SBURST, SRDY, SSIZE0, SSIZE1, SLOCK, SIRQ;

  buf  (RDATA0, SRDATA0);
  buf  (RDATA1, SRDATA1);
  buf  (RDATA2, SRDATA2);
  buf  (RDATA3, SRDATA3);
  buf  (RDATA4, SRDATA4);
  buf  (RDATA5, SRDATA5);
  buf  (RDATA6, SRDATA6);
  buf  (RDATA7, SRDATA7);
  buf  (RDATA8, SRDATA8);
  buf  (RDATA9, SRDATA9);
  buf  (RDATA10, SRDATA10);
  buf  (RDATA11, SRDATA11);
  buf  (RDATA12, SRDATA12);
  buf  (RDATA13, SRDATA13);
  buf  (RDATA14, SRDATA14);
  buf  (RDATA15, SRDATA15);
  buf  (RDATA16, SRDATA16);
  buf  (RDATA17, SRDATA17);
  buf  (RDATA18, SRDATA18);
  buf  (RDATA19, SRDATA19);
  buf  (RDATA20, SRDATA20);
  buf  (RDATA21, SRDATA21);
  buf  (RDATA22, SRDATA22);
  buf  (RDATA23, SRDATA23);
  buf  (RDATA24, SRDATA24);
  buf  (RDATA25, SRDATA25);
  buf  (RDATA26, SRDATA26);
  buf  (RDATA27, SRDATA27);
  buf  (RDATA28, SRDATA28);
  buf  (RDATA29, SRDATA29);
  buf  (RDATA30, SRDATA30);
  buf  (RDATA31, SRDATA31);
  buf  (RDATA32, SRDATA32);
  buf  (RDATA33, SRDATA33);
  buf  (RDATA34, SRDATA34);
  buf  (RDATA35, SRDATA35);
  buf  (GRANTED, SGRANTED);
  buf  (ACK, SACK);
  buf  (RETRY, SRETRY);
  buf  (ERR, SERR);
  buf  (SADDR0, ADDR0);
  buf  (SADDR1, ADDR1);
  buf  (SADDR2, ADDR2);
  buf  (SADDR3, ADDR3);
  buf  (SADDR4, ADDR4);
  buf  (SADDR5, ADDR5);
  buf  (SADDR6, ADDR6);
  buf  (SADDR7, ADDR7);
  buf  (SADDR8, ADDR8);
  buf  (SADDR9, ADDR9);
  buf  (SADDR10, ADDR10);
  buf  (SADDR11, ADDR11);
  buf  (SADDR12, ADDR12);
  buf  (SADDR13, ADDR13);
  buf  (SADDR14, ADDR14);
  buf  (SADDR15, ADDR15);
  buf  (SADDR16, ADDR16);
  buf  (SADDR17, ADDR17);
  buf  (SWDATA0, WDATA0);
  buf  (SWDATA1, WDATA1);
  buf  (SWDATA2, WDATA2);
  buf  (SWDATA3, WDATA3);
  buf  (SWDATA4, WDATA4);
  buf  (SWDATA5, WDATA5);
  buf  (SWDATA6, WDATA6);
  buf  (SWDATA7, WDATA7);
  buf  (SWDATA8, WDATA8);
  buf  (SWDATA9, WDATA9);
  buf  (SWDATA10, WDATA10);
  buf  (SWDATA11, WDATA11);
  buf  (SWDATA12, WDATA12);
  buf  (SWDATA13, WDATA13);
  buf  (SWDATA14, WDATA14);
  buf  (SWDATA15, WDATA15);
  buf  (SWDATA16, WDATA16);
  buf  (SWDATA17, WDATA17);
  buf  (SWDATA18, WDATA18);
  buf  (SWDATA19, WDATA19);
  buf  (SWDATA20, WDATA20);
  buf  (SWDATA21, WDATA21);
  buf  (SWDATA22, WDATA22);
  buf  (SWDATA23, WDATA23);
  buf  (SWDATA24, WDATA24);
  buf  (SWDATA25, WDATA25);
  buf  (SWDATA26, WDATA26);
  buf  (SWDATA27, WDATA27);
  buf  (SWDATA28, WDATA28);
  buf  (SWDATA29, WDATA29);
  buf  (SWDATA30, WDATA30);
  buf  (SWDATA31, WDATA31);
  buf  (SWDATA32, WDATA32);
  buf  (SWDATA33, WDATA33);
  buf  (SWDATA34, WDATA34);
  buf  (SWDATA35, WDATA35);
  buf  (SCLK, CLK);
  buf  (SRESET, RESET);
  buf  (SWRITE, WRITE);
  buf  (SREAD, READ);
  buf  (SBURST, BURST);
  buf  (SRDY, RDY);
  buf  (SSIZE0, SIZE0);
  buf  (SSIZE1, SIZE1);
  buf  (SLOCK, LOCK);
  buf  (SIRQ, IRQ);

endmodule

`endcelldefine

