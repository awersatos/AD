*Vacuum Tube Dual Triode (Audio freq.)
*Connections:
*              Plate 1
*              | Grid 1
*              | | Cathode 1
*              | | | Plate 2
*              | | | | Grid 2
*              | | | | | Cathode 2
*              | | | | | | H H
*              | | | | | | | |
.SUBCKT 6SN7   2 1 3 5 4 6 7 8
X1 2 1 3  6SN7s
X2 5 4 6 6SN7s
RH1 7 8 100
.ENDS 6SN7

*Vacuum Tube Triode (Audio freq.)
*Connections:
*            Plate
*            | Grid
*            | | Cathode
*            | | |
.SUBCKT 6SN7s 1 3 4
B1 2 4 I=((URAMP((V(2,4)/20)+V(3,4)))^1.5)/1086
C1 3 4 2.6E-12
C2 3 1 4.0E-12
C3 1 4 0.7E-12
R1 3 5 10E+3
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1.0E-12 RS=1.0)
.MODEL DX2 D(IS=1.0E-9 RS=1.0)
.ENDS 6SN7s
