*PIGBT
*P-IGBT Default  MCE  C G E  5-20-95
*MCE 600V 40A 24.3ns
*IGBT Pinout: 1=C, 2=G, 3=E
.SUBCKT PIGBT 71 72 74
Q1  83 81 85     QOUT
M1  81 82 83 83  MFIN L=1U W=1U
DSD 81 83  DO
DBE 81 85  DE
RC  85 71  21.2M
RE  83 73  2.12M
RG  72 82  25.5
CGE 82 83  1.42N
CGC 82 71  1P
EGD 91  0 81 82  1
VFB 93  0  0
FFB 81 82  VFB  1
CGD 92 93  1.41N
R1  92  0  1
D1  91 92  DLIM
DHV 94 93  DR
R2  91 94  1
D2  94  0  DLIM
LE  73 74  7.5N
DLV 94 95  DR 13
RLV 95  0  1
ESD 96 93  POLY(1) 81 83  19  1
MLV 95 96 93 93  SW
.MODEL SW NMOS (LEVEL=3 VTO=0 KP=5)
.MODEL QOUT NPN (IS=377F NF=1.2 BF=5.1 CJE=3.48N TF=24.3N XTB=1.3)
.MODEL MFIN PMOS (LEVEL=3 VMAX=400K THETA=46.1M ETA=2M VTO=-5.2 KP=2.12)
.MODEL DR D (IS=37.7F CJO=100P VJ=1 M=.82)
.MODEL DO D (IS=37.7F BV=600 CJO=2.07N VJ=1 M=.7)
.MODEL DE D (IS=37.7F BV=14.3 N=2)
.MODEL DLIM D (IS=100N)
.ENDS PIGBT
