*Vacuum Tube Pentode and Triode (Audio freq.)
*Connections:
*            Plate 1
*            | Grid 1
*            | | Cathode 1
*            | | | Plate 2
*            | | | | Grid 2
*            | | | | | Grid 3
*            | | | | | | Cathode 2
*            | | | | | | | Heater
*            | | | | | | | | Heater
*            | | | | | | | | |
.SUBCKT 7199 1 9 8 2 3 7 6 4 5
X1 1 9 8 7199T
X2 2 3 7 6 7199P
RH 4 5 100
.ENDS 7199

*Vacuum Tube Triode (Audio freq.)
*Connections:
*             Plate
*             | Grid
*             | | Cathode
*             | | |
.SUBCKT 7199T 1 3 4
B1 2 4 I=((URAMP((V(2,4)/17)+V(3,4)))^1.5)/711
C1 3 4 2.3E-12
C2 3 1 2.0E-12
C3 1 4 0.3E-12
R1 3 5 5E+3
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1.0E-12 RS=1.0)
.MODEL DX2 D(IS=1.0E-9 RS=1.0)
.ENDS 7199T

*Vacuum Tube Tetrode (Audio freq.)
*Connections:
*             Plate
*             | Screen
*             | | Grid
*             | | | Cathode
*             | | | |
.SUBCKT 7199P 1 6 3 4
B1 2 4 I=(((URAMP((V(7,4)/20)+V(3,4)))^1.5)/1206)*ATAN(V(1,4)/10)
B2 7 4 I=((URAMP((V(7,4)/20)+V(3,4)))^1.5)/2562
C1 3 4 5.0P
C2 3 1 0.06P
C3 1 4 2.0P
R1 3 5 5K
R2 2 4 2.5MEG
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
D4 6 7 DX
D5 4 7 DX2
.MODEL DX D(IS=1.0P RS=1.0)
.MODEL DX2 D(IS=1.0N RS=1.0)
.ENDS 7199P